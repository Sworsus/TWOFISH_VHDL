----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:40:58 04/21/2021 
-- Design Name: 
-- Module Name:    mult_EF_mem - mult_EF_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mult_EF_mem is
	port (
			in_EF : in STD_LOGIC_VECTOR (7 downto 0);
			out_EF : out STD_LOGIC_VECTOR (7 downto 0)
			);	
end mult_EF_mem;

architecture mult_EF_mem of mult_EF_mem is
begin
	with in_EF select
		out_EF <=	"00000000" when "00000000", "11101111" when "00000001", "10110111" when "00000010", "01011000" when "00000011", 
						"00000111" when "00000100", "11101000" when "00000101", "10110000" when "00000110", "01011111" when "00000111", 
						"00001110" when "00001000", "11100001" when "00001001", "10111001" when "00001010", "01010110" when "00001011", 
						"00001001" when "00001100", "11100110" when "00001101", "10111110" when "00001110", "01010001" when "00001111", 
						"00011100" when "00010000", "11110011" when "00010001", "10101011" when "00010010", "01000100" when "00010011", 
						"00011011" when "00010100", "11110100" when "00010101", "10101100" when "00010110", "01000011" when "00010111", 
						"00010010" when "00011000", "11111101" when "00011001", "10100101" when "00011010", "01001010" when "00011011", 
						"00010101" when "00011100", "11111010" when "00011101", "10100010" when "00011110", "01001101" when "00011111", 
						"00111000" when "00100000", "11010111" when "00100001", "10001111" when "00100010", "01100000" when "00100011", 
						"00111111" when "00100100", "11010000" when "00100101", "10001000" when "00100110", "01100111" when "00100111", 
						"00110110" when "00101000", "11011001" when "00101001", "10000001" when "00101010", "01101110" when "00101011", 
						"00110001" when "00101100", "11011110" when "00101101", "10000110" when "00101110", "01101001" when "00101111", 
						"00100100" when "00110000", "11001011" when "00110001", "10010011" when "00110010", "01111100" when "00110011", 
						"00100011" when "00110100", "11001100" when "00110101", "10010100" when "00110110", "01111011" when "00110111", 
						"00101010" when "00111000", "11000101" when "00111001", "10011101" when "00111010", "01110010" when "00111011", 
						"00101101" when "00111100", "11000010" when "00111101", "10011010" when "00111110", "01110101" when "00111111", 
						"01110000" when "01000000", "10011111" when "01000001", "11000111" when "01000010", "00101000" when "01000011", 
						"01110111" when "01000100", "10011000" when "01000101", "11000000" when "01000110", "00101111" when "01000111", 
						"01111110" when "01001000", "10010001" when "01001001", "11001001" when "01001010", "00100110" when "01001011", 
						"01111001" when "01001100", "10010110" when "01001101", "11001110" when "01001110", "00100001" when "01001111", 
						"01101100" when "01010000", "10000011" when "01010001", "11011011" when "01010010", "00110100" when "01010011", 
						"01101011" when "01010100", "10000100" when "01010101", "11011100" when "01010110", "00110011" when "01010111", 
						"01100010" when "01011000", "10001101" when "01011001", "11010101" when "01011010", "00111010" when "01011011", 
						"01100101" when "01011100", "10001010" when "01011101", "11010010" when "01011110", "00111101" when "01011111", 
						"01001000" when "01100000", "10100111" when "01100001", "11111111" when "01100010", "00010000" when "01100011", 
						"01001111" when "01100100", "10100000" when "01100101", "11111000" when "01100110", "00010111" when "01100111", 
						"01000110" when "01101000", "10101001" when "01101001", "11110001" when "01101010", "00011110" when "01101011", 
						"01000001" when "01101100", "10101110" when "01101101", "11110110" when "01101110", "00011001" when "01101111", 
						"01010100" when "01110000", "10111011" when "01110001", "11100011" when "01110010", "00001100" when "01110011", 
						"01010011" when "01110100", "10111100" when "01110101", "11100100" when "01110110", "00001011" when "01110111", 
						"01011010" when "01111000", "10110101" when "01111001", "11101101" when "01111010", "00000010" when "01111011", 
						"01011101" when "01111100", "10110010" when "01111101", "11101010" when "01111110", "00000101" when "01111111", 
						"11100000" when "10000000", "00001111" when "10000001", "01010111" when "10000010", "10111000" when "10000011", 
						"11100111" when "10000100", "00001000" when "10000101", "01010000" when "10000110", "10111111" when "10000111", 
						"11101110" when "10001000", "00000001" when "10001001", "01011001" when "10001010", "10110110" when "10001011", 
						"11101001" when "10001100", "00000110" when "10001101", "01011110" when "10001110", "10110001" when "10001111", 
						"11111100" when "10010000", "00010011" when "10010001", "01001011" when "10010010", "10100100" when "10010011", 
						"11111011" when "10010100", "00010100" when "10010101", "01001100" when "10010110", "10100011" when "10010111", 
						"11110010" when "10011000", "00011101" when "10011001", "01000101" when "10011010", "10101010" when "10011011", 
						"11110101" when "10011100", "00011010" when "10011101", "01000010" when "10011110", "10101101" when "10011111", 
						"11011000" when "10100000", "00110111" when "10100001", "01101111" when "10100010", "10000000" when "10100011", 
						"11011111" when "10100100", "00110000" when "10100101", "01101000" when "10100110", "10000111" when "10100111", 
						"11010110" when "10101000", "00111001" when "10101001", "01100001" when "10101010", "10001110" when "10101011", 
						"11010001" when "10101100", "00111110" when "10101101", "01100110" when "10101110", "10001001" when "10101111", 
						"11000100" when "10110000", "00101011" when "10110001", "01110011" when "10110010", "10011100" when "10110011", 
						"11000011" when "10110100", "00101100" when "10110101", "01110100" when "10110110", "10011011" when "10110111", 
						"11001010" when "10111000", "00100101" when "10111001", "01111101" when "10111010", "10010010" when "10111011", 
						"11001101" when "10111100", "00100010" when "10111101", "01111010" when "10111110", "10010101" when "10111111", 
						"10010000" when "11000000", "01111111" when "11000001", "00100111" when "11000010", "11001000" when "11000011", 
						"10010111" when "11000100", "01111000" when "11000101", "00100000" when "11000110", "11001111" when "11000111", 
						"10011110" when "11001000", "01110001" when "11001001", "00101001" when "11001010", "11000110" when "11001011", 
						"10011001" when "11001100", "01110110" when "11001101", "00101110" when "11001110", "11000001" when "11001111", 
						"10001100" when "11010000", "01100011" when "11010001", "00111011" when "11010010", "11010100" when "11010011", 
						"10001011" when "11010100", "01100100" when "11010101", "00111100" when "11010110", "11010011" when "11010111", 
						"10000010" when "11011000", "01101101" when "11011001", "00110101" when "11011010", "11011010" when "11011011", 
						"10000101" when "11011100", "01101010" when "11011101", "00110010" when "11011110", "11011101" when "11011111", 
						"10101000" when "11100000", "01000111" when "11100001", "00011111" when "11100010", "11110000" when "11100011", 
						"10101111" when "11100100", "01000000" when "11100101", "00011000" when "11100110", "11110111" when "11100111", 
						"10100110" when "11101000", "01001001" when "11101001", "00010001" when "11101010", "11111110" when "11101011", 
						"10100001" when "11101100", "01001110" when "11101101", "00010110" when "11101110", "11111001" when "11101111", 
						"10110100" when "11110000", "01011011" when "11110001", "00000011" when "11110010", "11101100" when "11110011", 
						"10110011" when "11110100", "01011100" when "11110101", "00000100" when "11110110", "11101011" when "11110111", 
						"10111010" when "11111000", "01010101" when "11111001", "00001101" when "11111010", "11100010" when "11111011", 
						"10111101" when "11111100", "01010010" when "11111101", "00001010" when "11111110", "11100101" when "11111111";
end mult_EF_mem;

