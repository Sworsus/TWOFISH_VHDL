----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    00:41:43 04/24/2021 
-- Design Name: 
-- Module Name:    mul_47_mem - mul_47_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_47_mem is
	port (
			in_47 : in STD_LOGIC_VECTOR (7 downto 0);
			out_47 : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_47_mem;

architecture mul_47_mem of mul_47_mem is
begin
	with in_47 select
		out_47 <= "00000000" when "00000000", 
					"01000111" when "00000001", 
					"10001110" when "00000010", 
					"11001001" when "00000011", 
					"01110101" when "00000100", 
					"00110010" when "00000101", 
					"11111011" when "00000110", 
					"10111100" when "00000111", 
					"11101010" when "00001000", 
					"10101101" when "00001001", 
					"01100100" when "00001010", 
					"00100011" when "00001011", 
					"10011111" when "00001100", 
					"11011000" when "00001101", 
					"00010001" when "00001110", 
					"01010110" when "00001111", 
					"10111101" when "00010000", 
					"11111010" when "00010001", 
					"00110011" when "00010010", 
					"01110100" when "00010011", 
					"11001000" when "00010100", 
					"10001111" when "00010101", 
					"01000110" when "00010110", 
					"00000001" when "00010111", 
					"01010111" when "00011000", 
					"00010000" when "00011001", 
					"11011001" when "00011010", 
					"10011110" when "00011011", 
					"00100010" when "00011100", 
					"01100101" when "00011101", 
					"10101100" when "00011110", 
					"11101011" when "00011111", 
					"00010011" when "00100000", 
					"01010100" when "00100001", 
					"10011101" when "00100010", 
					"11011010" when "00100011", 
					"01100110" when "00100100", 
					"00100001" when "00100101", 
					"11101000" when "00100110", 
					"10101111" when "00100111", 
					"11111001" when "00101000", 
					"10111110" when "00101001", 
					"01110111" when "00101010", 
					"00110000" when "00101011", 
					"10001100" when "00101100", 
					"11001011" when "00101101", 
					"00000010" when "00101110", 
					"01000101" when "00101111", 
					"10101110" when "00110000", 
					"11101001" when "00110001", 
					"00100000" when "00110010", 
					"01100111" when "00110011", 
					"11011011" when "00110100", 
					"10011100" when "00110101", 
					"01010101" when "00110110", 
					"00010010" when "00110111", 
					"01000100" when "00111000", 
					"00000011" when "00111001", 
					"11001010" when "00111010", 
					"10001101" when "00111011", 
					"00110001" when "00111100", 
					"01110110" when "00111101", 
					"10111111" when "00111110", 
					"11111000" when "00111111", 
					"00100110" when "01000000", 
					"01100001" when "01000001", 
					"10101000" when "01000010", 
					"11101111" when "01000011", 
					"01010011" when "01000100", 
					"00010100" when "01000101", 
					"11011101" when "01000110", 
					"10011010" when "01000111", 
					"11001100" when "01001000", 
					"10001011" when "01001001", 
					"01000010" when "01001010", 
					"00000101" when "01001011", 
					"10111001" when "01001100", 
					"11111110" when "01001101", 
					"00110111" when "01001110", 
					"01110000" when "01001111", 
					"10011011" when "01010000", 
					"11011100" when "01010001", 
					"00010101" when "01010010", 
					"01010010" when "01010011", 
					"11101110" when "01010100", 
					"10101001" when "01010101", 
					"01100000" when "01010110", 
					"00100111" when "01010111", 
					"01110001" when "01011000", 
					"00110110" when "01011001", 
					"11111111" when "01011010", 
					"10111000" when "01011011", 
					"00000100" when "01011100", 
					"01000011" when "01011101", 
					"10001010" when "01011110", 
					"11001101" when "01011111", 
					"00110101" when "01100000", 
					"01110010" when "01100001", 
					"10111011" when "01100010", 
					"11111100" when "01100011", 
					"01000000" when "01100100", 
					"00000111" when "01100101", 
					"11001110" when "01100110", 
					"10001001" when "01100111", 
					"11011111" when "01101000", 
					"10011000" when "01101001", 
					"01010001" when "01101010", 
					"00010110" when "01101011", 
					"10101010" when "01101100", 
					"11101101" when "01101101", 
					"00100100" when "01101110", 
					"01100011" when "01101111", 
					"10001000" when "01110000", 
					"11001111" when "01110001", 
					"00000110" when "01110010", 
					"01000001" when "01110011", 
					"11111101" when "01110100", 
					"10111010" when "01110101", 
					"01110011" when "01110110", 
					"00110100" when "01110111", 
					"01100010" when "01111000", 
					"00100101" when "01111001", 
					"11101100" when "01111010", 
					"10101011" when "01111011", 
					"00010111" when "01111100", 
					"01010000" when "01111101", 
					"10011001" when "01111110", 
					"11011110" when "01111111", 
					"01001100" when "10000000", 
					"00001011" when "10000001", 
					"11000010" when "10000010", 
					"10000101" when "10000011", 
					"00111001" when "10000100", 
					"01111110" when "10000101", 
					"10110111" when "10000110", 
					"11110000" when "10000111", 
					"10100110" when "10001000", 
					"11100001" when "10001001", 
					"00101000" when "10001010", 
					"01101111" when "10001011", 
					"11010011" when "10001100", 
					"10010100" when "10001101", 
					"01011101" when "10001110", 
					"00011010" when "10001111", 
					"11110001" when "10010000", 
					"10110110" when "10010001", 
					"01111111" when "10010010", 
					"00111000" when "10010011", 
					"10000100" when "10010100", 
					"11000011" when "10010101", 
					"00001010" when "10010110", 
					"01001101" when "10010111", 
					"00011011" when "10011000", 
					"01011100" when "10011001", 
					"10010101" when "10011010", 
					"11010010" when "10011011", 
					"01101110" when "10011100", 
					"00101001" when "10011101", 
					"11100000" when "10011110", 
					"10100111" when "10011111", 
					"01011111" when "10100000", 
					"00011000" when "10100001", 
					"11010001" when "10100010", 
					"10010110" when "10100011", 
					"00101010" when "10100100", 
					"01101101" when "10100101", 
					"10100100" when "10100110", 
					"11100011" when "10100111", 
					"10110101" when "10101000", 
					"11110010" when "10101001", 
					"00111011" when "10101010", 
					"01111100" when "10101011", 
					"11000000" when "10101100", 
					"10000111" when "10101101", 
					"01001110" when "10101110", 
					"00001001" when "10101111", 
					"11100010" when "10110000", 
					"10100101" when "10110001", 
					"01101100" when "10110010", 
					"00101011" when "10110011", 
					"10010111" when "10110100", 
					"11010000" when "10110101", 
					"00011001" when "10110110", 
					"01011110" when "10110111", 
					"00001000" when "10111000", 
					"01001111" when "10111001", 
					"10000110" when "10111010", 
					"11000001" when "10111011", 
					"01111101" when "10111100", 
					"00111010" when "10111101", 
					"11110011" when "10111110", 
					"10110100" when "10111111", 
					"01101010" when "11000000", 
					"00101101" when "11000001", 
					"11100100" when "11000010", 
					"10100011" when "11000011", 
					"00011111" when "11000100", 
					"01011000" when "11000101", 
					"10010001" when "11000110", 
					"11010110" when "11000111", 
					"10000000" when "11001000", 
					"11000111" when "11001001", 
					"00001110" when "11001010", 
					"01001001" when "11001011", 
					"11110101" when "11001100", 
					"10110010" when "11001101", 
					"01111011" when "11001110", 
					"00111100" when "11001111", 
					"11010111" when "11010000", 
					"10010000" when "11010001", 
					"01011001" when "11010010", 
					"00011110" when "11010011", 
					"10100010" when "11010100", 
					"11100101" when "11010101", 
					"00101100" when "11010110", 
					"01101011" when "11010111", 
					"00111101" when "11011000", 
					"01111010" when "11011001", 
					"10110011" when "11011010", 
					"11110100" when "11011011", 
					"01001000" when "11011100", 
					"00001111" when "11011101", 
					"11000110" when "11011110", 
					"10000001" when "11011111", 
					"01111001" when "11100000", 
					"00111110" when "11100001", 
					"11110111" when "11100010", 
					"10110000" when "11100011", 
					"00001100" when "11100100", 
					"01001011" when "11100101", 
					"10000010" when "11100110", 
					"11000101" when "11100111", 
					"10010011" when "11101000", 
					"11010100" when "11101001", 
					"00011101" when "11101010", 
					"01011010" when "11101011", 
					"11100110" when "11101100", 
					"10100001" when "11101101", 
					"01101000" when "11101110", 
					"00101111" when "11101111", 
					"11000100" when "11110000", 
					"10000011" when "11110001", 
					"01001010" when "11110010", 
					"00001101" when "11110011", 
					"10110001" when "11110100", 
					"11110110" when "11110101", 
					"00111111" when "11110110", 
					"01111000" when "11110111", 
					"00101110" when "11111000", 
					"01101001" when "11111001", 
					"10100000" when "11111010", 
					"11100111" when "11111011", 
					"01011011" when "11111100", 
					"00011100" when "11111101", 
					"11010101" when "11111110", 
					"10010010" when "11111111";

end mul_47_mem;

