----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:39:15 04/24/2021 
-- Design Name: 
-- Module Name:    mul_87_mem - mul_87_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_87_mem is
	port (
			in_87 : in STD_LOGIC_VECTOR (7 downto 0);
			out_87 : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_87_mem;

architecture mul_87_mem of mul_87_mem is

begin

	with in_87 select
	out_87 <= "00000000" when "00000000", 
				"10000111" when "00000001", 
				"01100111" when "00000010", 
				"11100000" when "00000011", 
				"11001110" when "00000100", 
				"01001001" when "00000101", 
				"10101001" when "00000110", 
				"00101110" when "00000111", 
				"11110101" when "00001000", 
				"01110010" when "00001001", 
				"10010010" when "00001010", 
				"00010101" when "00001011", 
				"00111011" when "00001100", 
				"10111100" when "00001101", 
				"01011100" when "00001110", 
				"11011011" when "00001111", 
				"10000011" when "00010000", 
				"00000100" when "00010001", 
				"11100100" when "00010010", 
				"01100011" when "00010011", 
				"01001101" when "00010100", 
				"11001010" when "00010101", 
				"00101010" when "00010110", 
				"10101101" when "00010111", 
				"01110110" when "00011000", 
				"11110001" when "00011001", 
				"00010001" when "00011010", 
				"10010110" when "00011011", 
				"10111000" when "00011100", 
				"00111111" when "00011101", 
				"11011111" when "00011110", 
				"01011000" when "00011111", 
				"01101111" when "00100000", 
				"11101000" when "00100001", 
				"00001000" when "00100010", 
				"10001111" when "00100011", 
				"10100001" when "00100100", 
				"00100110" when "00100101", 
				"11000110" when "00100110", 
				"01000001" when "00100111", 
				"10011010" when "00101000", 
				"00011101" when "00101001", 
				"11111101" when "00101010", 
				"01111010" when "00101011", 
				"01010100" when "00101100", 
				"11010011" when "00101101", 
				"00110011" when "00101110", 
				"10110100" when "00101111", 
				"11101100" when "00110000", 
				"01101011" when "00110001", 
				"10001011" when "00110010", 
				"00001100" when "00110011", 
				"00100010" when "00110100", 
				"10100101" when "00110101", 
				"01000101" when "00110110", 
				"11000010" when "00110111", 
				"00011001" when "00111000", 
				"10011110" when "00111001", 
				"01111110" when "00111010", 
				"11111001" when "00111011", 
				"11010111" when "00111100", 
				"01010000" when "00111101", 
				"10110000" when "00111110", 
				"00110111" when "00111111", 
				"11011110" when "01000000", 
				"01011001" when "01000001", 
				"10111001" when "01000010", 
				"00111110" when "01000011", 
				"00010000" when "01000100", 
				"10010111" when "01000101", 
				"01110111" when "01000110", 
				"11110000" when "01000111", 
				"00101011" when "01001000", 
				"10101100" when "01001001", 
				"01001100" when "01001010", 
				"11001011" when "01001011", 
				"11100101" when "01001100", 
				"01100010" when "01001101", 
				"10000010" when "01001110", 
				"00000101" when "01001111", 
				"01011101" when "01010000", 
				"11011010" when "01010001", 
				"00111010" when "01010010", 
				"10111101" when "01010011", 
				"10010011" when "01010100", 
				"00010100" when "01010101", 
				"11110100" when "01010110", 
				"01110011" when "01010111", 
				"10101000" when "01011000", 
				"00101111" when "01011001", 
				"11001111" when "01011010", 
				"01001000" when "01011011", 
				"01100110" when "01011100", 
				"11100001" when "01011101", 
				"00000001" when "01011110", 
				"10000110" when "01011111", 
				"10110001" when "01100000", 
				"00110110" when "01100001", 
				"11010110" when "01100010", 
				"01010001" when "01100011", 
				"01111111" when "01100100", 
				"11111000" when "01100101", 
				"00011000" when "01100110", 
				"10011111" when "01100111", 
				"01000100" when "01101000", 
				"11000011" when "01101001", 
				"00100011" when "01101010", 
				"10100100" when "01101011", 
				"10001010" when "01101100", 
				"00001101" when "01101101", 
				"11101101" when "01101110", 
				"01101010" when "01101111", 
				"00110010" when "01110000", 
				"10110101" when "01110001", 
				"01010101" when "01110010", 
				"11010010" when "01110011", 
				"11111100" when "01110100", 
				"01111011" when "01110101", 
				"10011011" when "01110110", 
				"00011100" when "01110111", 
				"11000111" when "01111000", 
				"01000000" when "01111001", 
				"10100000" when "01111010", 
				"00100111" when "01111011", 
				"00001001" when "01111100", 
				"10001110" when "01111101", 
				"01101110" when "01111110", 
				"11101001" when "01111111", 
				"11010101" when "10000000", 
				"01010010" when "10000001", 
				"10110010" when "10000010", 
				"00110101" when "10000011", 
				"00011011" when "10000100", 
				"10011100" when "10000101", 
				"01111100" when "10000110", 
				"11111011" when "10000111", 
				"00100000" when "10001000", 
				"10100111" when "10001001", 
				"01000111" when "10001010", 
				"11000000" when "10001011", 
				"11101110" when "10001100", 
				"01101001" when "10001101", 
				"10001001" when "10001110", 
				"00001110" when "10001111", 
				"01010110" when "10010000", 
				"11010001" when "10010001", 
				"00110001" when "10010010", 
				"10110110" when "10010011", 
				"10011000" when "10010100", 
				"00011111" when "10010101", 
				"11111111" when "10010110", 
				"01111000" when "10010111", 
				"10100011" when "10011000", 
				"00100100" when "10011001", 
				"11000100" when "10011010", 
				"01000011" when "10011011", 
				"01101101" when "10011100", 
				"11101010" when "10011101", 
				"00001010" when "10011110", 
				"10001101" when "10011111", 
				"10111010" when "10100000", 
				"00111101" when "10100001", 
				"11011101" when "10100010", 
				"01011010" when "10100011", 
				"01110100" when "10100100", 
				"11110011" when "10100101", 
				"00010011" when "10100110", 
				"10010100" when "10100111", 
				"01001111" when "10101000", 
				"11001000" when "10101001", 
				"00101000" when "10101010", 
				"10101111" when "10101011", 
				"10000001" when "10101100", 
				"00000110" when "10101101", 
				"11100110" when "10101110", 
				"01100001" when "10101111", 
				"00111001" when "10110000", 
				"10111110" when "10110001", 
				"01011110" when "10110010", 
				"11011001" when "10110011", 
				"11110111" when "10110100", 
				"01110000" when "10110101", 
				"10010000" when "10110110", 
				"00010111" when "10110111", 
				"11001100" when "10111000", 
				"01001011" when "10111001", 
				"10101011" when "10111010", 
				"00101100" when "10111011", 
				"00000010" when "10111100", 
				"10000101" when "10111101", 
				"01100101" when "10111110", 
				"11100010" when "10111111", 
				"00001011" when "11000000", 
				"10001100" when "11000001", 
				"01101100" when "11000010", 
				"11101011" when "11000011", 
				"11000101" when "11000100", 
				"01000010" when "11000101", 
				"10100010" when "11000110", 
				"00100101" when "11000111", 
				"11111110" when "11001000", 
				"01111001" when "11001001", 
				"10011001" when "11001010", 
				"00011110" when "11001011", 
				"00110000" when "11001100", 
				"10110111" when "11001101", 
				"01010111" when "11001110", 
				"11010000" when "11001111", 
				"10001000" when "11010000", 
				"00001111" when "11010001", 
				"11101111" when "11010010", 
				"01101000" when "11010011", 
				"01000110" when "11010100", 
				"11000001" when "11010101", 
				"00100001" when "11010110", 
				"10100110" when "11010111", 
				"01111101" when "11011000", 
				"11111010" when "11011001", 
				"00011010" when "11011010", 
				"10011101" when "11011011", 
				"10110011" when "11011100", 
				"00110100" when "11011101", 
				"11010100" when "11011110", 
				"01010011" when "11011111", 
				"01100100" when "11100000", 
				"11100011" when "11100001", 
				"00000011" when "11100010", 
				"10000100" when "11100011", 
				"10101010" when "11100100", 
				"00101101" when "11100101", 
				"11001101" when "11100110", 
				"01001010" when "11100111", 
				"10010001" when "11101000", 
				"00010110" when "11101001", 
				"11110110" when "11101010", 
				"01110001" when "11101011", 
				"01011111" when "11101100", 
				"11011000" when "11101101", 
				"00111000" when "11101110", 
				"10111111" when "11101111", 
				"11100111" when "11110000", 
				"01100000" when "11110001", 
				"10000000" when "11110010", 
				"00000111" when "11110011", 
				"00101001" when "11110100", 
				"10101110" when "11110101", 
				"01001110" when "11110110", 
				"11001001" when "11110111", 
				"00010010" when "11111000", 
				"10010101" when "11111001", 
				"01110101" when "11111010", 
				"11110010" when "11111011", 
				"11011100" when "11111100", 
				"01011011" when "11111101", 
				"10111011" when "11111110", 
				"00111100" when "11111111";

end mul_87_mem;

