----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:37:57 04/24/2021 
-- Design Name: 
-- Module Name:    mul_C1_mem - mul_C1_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_C1_mem is
	port (
			in_C1 : in STD_LOGIC_VECTOR (7 downto 0);
			out_C1 : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_C1_mem;

architecture mul_C1_mem of mul_C1_mem is

begin

	with in_C1 select
	out_C1 <= "00000000" when "00000000", 
				"11000001" when "00000001", 
				"11101011" when "00000010", 
				"00101010" when "00000011", 
				"10111111" when "00000100", 
				"01111110" when "00000101", 
				"01010100" when "00000110", 
				"10010101" when "00000111", 
				"00010111" when "00001000", 
				"11010110" when "00001001", 
				"11111100" when "00001010", 
				"00111101" when "00001011", 
				"10101000" when "00001100", 
				"01101001" when "00001101", 
				"01000011" when "00001110", 
				"10000010" when "00001111", 
				"00101110" when "00010000", 
				"11101111" when "00010001", 
				"11000101" when "00010010", 
				"00000100" when "00010011", 
				"10010001" when "00010100", 
				"01010000" when "00010101", 
				"01111010" when "00010110", 
				"10111011" when "00010111", 
				"00111001" when "00011000", 
				"11111000" when "00011001", 
				"11010010" when "00011010", 
				"00010011" when "00011011", 
				"10000110" when "00011100", 
				"01000111" when "00011101", 
				"01101101" when "00011110", 
				"10101100" when "00011111", 
				"01011100" when "00100000", 
				"10011101" when "00100001", 
				"10110111" when "00100010", 
				"01110110" when "00100011", 
				"11100011" when "00100100", 
				"00100010" when "00100101", 
				"00001000" when "00100110", 
				"11001001" when "00100111", 
				"01001011" when "00101000", 
				"10001010" when "00101001", 
				"10100000" when "00101010", 
				"01100001" when "00101011", 
				"11110100" when "00101100", 
				"00110101" when "00101101", 
				"00011111" when "00101110", 
				"11011110" when "00101111", 
				"01110010" when "00110000", 
				"10110011" when "00110001", 
				"10011001" when "00110010", 
				"01011000" when "00110011", 
				"11001101" when "00110100", 
				"00001100" when "00110101", 
				"00100110" when "00110110", 
				"11100111" when "00110111", 
				"01100101" when "00111000", 
				"10100100" when "00111001", 
				"10001110" when "00111010", 
				"01001111" when "00111011", 
				"11011010" when "00111100", 
				"00011011" when "00111101", 
				"00110001" when "00111110", 
				"11110000" when "00111111", 
				"10111000" when "01000000", 
				"01111001" when "01000001", 
				"01010011" when "01000010", 
				"10010010" when "01000011", 
				"00000111" when "01000100", 
				"11000110" when "01000101", 
				"11101100" when "01000110", 
				"00101101" when "01000111", 
				"10101111" when "01001000", 
				"01101110" when "01001001", 
				"01000100" when "01001010", 
				"10000101" when "01001011", 
				"00010000" when "01001100", 
				"11010001" when "01001101", 
				"11111011" when "01001110", 
				"00111010" when "01001111", 
				"10010110" when "01010000", 
				"01010111" when "01010001", 
				"01111101" when "01010010", 
				"10111100" when "01010011", 
				"00101001" when "01010100", 
				"11101000" when "01010101", 
				"11000010" when "01010110", 
				"00000011" when "01010111", 
				"10000001" when "01011000", 
				"01000000" when "01011001", 
				"01101010" when "01011010", 
				"10101011" when "01011011", 
				"00111110" when "01011100", 
				"11111111" when "01011101", 
				"11010101" when "01011110", 
				"00010100" when "01011111", 
				"11100100" when "01100000", 
				"00100101" when "01100001", 
				"00001111" when "01100010", 
				"11001110" when "01100011", 
				"01011011" when "01100100", 
				"10011010" when "01100101", 
				"10110000" when "01100110", 
				"01110001" when "01100111", 
				"11110011" when "01101000", 
				"00110010" when "01101001", 
				"00011000" when "01101010", 
				"11011001" when "01101011", 
				"01001100" when "01101100", 
				"10001101" when "01101101", 
				"10100111" when "01101110", 
				"01100110" when "01101111", 
				"11001010" when "01110000", 
				"00001011" when "01110001", 
				"00100001" when "01110010", 
				"11100000" when "01110011", 
				"01110101" when "01110100", 
				"10110100" when "01110101", 
				"10011110" when "01110110", 
				"01011111" when "01110111", 
				"11011101" when "01111000", 
				"00011100" when "01111001", 
				"00110110" when "01111010", 
				"11110111" when "01111011", 
				"01100010" when "01111100", 
				"10100011" when "01111101", 
				"10001001" when "01111110", 
				"01001000" when "01111111", 
				"00011001" when "10000000", 
				"11011000" when "10000001", 
				"11110010" when "10000010", 
				"00110011" when "10000011", 
				"10100110" when "10000100", 
				"01100111" when "10000101", 
				"01001101" when "10000110", 
				"10001100" when "10000111", 
				"00001110" when "10001000", 
				"11001111" when "10001001", 
				"11100101" when "10001010", 
				"00100100" when "10001011", 
				"10110001" when "10001100", 
				"01110000" when "10001101", 
				"01011010" when "10001110", 
				"10011011" when "10001111", 
				"00110111" when "10010000", 
				"11110110" when "10010001", 
				"11011100" when "10010010", 
				"00011101" when "10010011", 
				"10001000" when "10010100", 
				"01001001" when "10010101", 
				"01100011" when "10010110", 
				"10100010" when "10010111", 
				"00100000" when "10011000", 
				"11100001" when "10011001", 
				"11001011" when "10011010", 
				"00001010" when "10011011", 
				"10011111" when "10011100", 
				"01011110" when "10011101", 
				"01110100" when "10011110", 
				"10110101" when "10011111", 
				"01000101" when "10100000", 
				"10000100" when "10100001", 
				"10101110" when "10100010", 
				"01101111" when "10100011", 
				"11111010" when "10100100", 
				"00111011" when "10100101", 
				"00010001" when "10100110", 
				"11010000" when "10100111", 
				"01010010" when "10101000", 
				"10010011" when "10101001", 
				"10111001" when "10101010", 
				"01111000" when "10101011", 
				"11101101" when "10101100", 
				"00101100" when "10101101", 
				"00000110" when "10101110", 
				"11000111" when "10101111", 
				"01101011" when "10110000", 
				"10101010" when "10110001", 
				"10000000" when "10110010", 
				"01000001" when "10110011", 
				"11010100" when "10110100", 
				"00010101" when "10110101", 
				"00111111" when "10110110", 
				"11111110" when "10110111", 
				"01111100" when "10111000", 
				"10111101" when "10111001", 
				"10010111" when "10111010", 
				"01010110" when "10111011", 
				"11000011" when "10111100", 
				"00000010" when "10111101", 
				"00101000" when "10111110", 
				"11101001" when "10111111", 
				"10100001" when "11000000", 
				"01100000" when "11000001", 
				"01001010" when "11000010", 
				"10001011" when "11000011", 
				"00011110" when "11000100", 
				"11011111" when "11000101", 
				"11110101" when "11000110", 
				"00110100" when "11000111", 
				"10110110" when "11001000", 
				"01110111" when "11001001", 
				"01011101" when "11001010", 
				"10011100" when "11001011", 
				"00001001" when "11001100", 
				"11001000" when "11001101", 
				"11100010" when "11001110", 
				"00100011" when "11001111", 
				"10001111" when "11010000", 
				"01001110" when "11010001", 
				"01100100" when "11010010", 
				"10100101" when "11010011", 
				"00110000" when "11010100", 
				"11110001" when "11010101", 
				"11011011" when "11010110", 
				"00011010" when "11010111", 
				"10011000" when "11011000", 
				"01011001" when "11011001", 
				"01110011" when "11011010", 
				"10110010" when "11011011", 
				"00100111" when "11011100", 
				"11100110" when "11011101", 
				"11001100" when "11011110", 
				"00001101" when "11011111", 
				"11111101" when "11100000", 
				"00111100" when "11100001", 
				"00010110" when "11100010", 
				"11010111" when "11100011", 
				"01000010" when "11100100", 
				"10000011" when "11100101", 
				"10101001" when "11100110", 
				"01101000" when "11100111", 
				"11101010" when "11101000", 
				"00101011" when "11101001", 
				"00000001" when "11101010", 
				"11000000" when "11101011", 
				"01010101" when "11101100", 
				"10010100" when "11101101", 
				"10111110" when "11101110", 
				"01111111" when "11101111", 
				"11010011" when "11110000", 
				"00010010" when "11110001", 
				"00111000" when "11110010", 
				"11111001" when "11110011", 
				"01101100" when "11110100", 
				"10101101" when "11110101", 
				"10000111" when "11110110", 
				"01000110" when "11110111", 
				"11000100" when "11111000", 
				"00000101" when "11111001", 
				"00101111" when "11111010", 
				"11101110" when "11111011", 
				"01111011" when "11111100", 
				"10111010" when "11111101", 
				"10010000" when "11111110", 
				"01010001" when "11111111";

end mul_C1_mem;

