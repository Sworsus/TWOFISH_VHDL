----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:01:36 04/24/2021 
-- Design Name: 
-- Module Name:    mul_E5_mem - mul_E5_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_E5_mem is
	port (
			in_E5 : in STD_LOGIC_VECTOR (7 downto 0);
			out_E5 : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_E5_mem;

architecture mul_E5_mem of mul_E5_mem is

begin

	with in_E5 select
	out_E5 <= "00000000" when "00000000", 
				"11100101" when "00000001", 
				"10100011" when "00000010", 
				"01000110" when "00000011", 
				"00101111" when "00000100", 
				"11001010" when "00000101", 
				"10001100" when "00000110", 
				"01101001" when "00000111", 
				"01011110" when "00001000", 
				"10111011" when "00001001", 
				"11111101" when "00001010", 
				"00011000" when "00001011", 
				"01110001" when "00001100", 
				"10010100" when "00001101", 
				"11010010" when "00001110", 
				"00110111" when "00001111", 
				"10111100" when "00010000", 
				"01011001" when "00010001", 
				"00011111" when "00010010", 
				"11111010" when "00010011", 
				"10010011" when "00010100", 
				"01110110" when "00010101", 
				"00110000" when "00010110", 
				"11010101" when "00010111", 
				"11100010" when "00011000", 
				"00000111" when "00011001", 
				"01000001" when "00011010", 
				"10100100" when "00011011", 
				"11001101" when "00011100", 
				"00101000" when "00011101", 
				"01101110" when "00011110", 
				"10001011" when "00011111", 
				"00010001" when "00100000", 
				"11110100" when "00100001", 
				"10110010" when "00100010", 
				"01010111" when "00100011", 
				"00111110" when "00100100", 
				"11011011" when "00100101", 
				"10011101" when "00100110", 
				"01111000" when "00100111", 
				"01001111" when "00101000", 
				"10101010" when "00101001", 
				"11101100" when "00101010", 
				"00001001" when "00101011", 
				"01100000" when "00101100", 
				"10000101" when "00101101", 
				"11000011" when "00101110", 
				"00100110" when "00101111", 
				"10101101" when "00110000", 
				"01001000" when "00110001", 
				"00001110" when "00110010", 
				"11101011" when "00110011", 
				"10000010" when "00110100", 
				"01100111" when "00110101", 
				"00100001" when "00110110", 
				"11000100" when "00110111", 
				"11110011" when "00111000", 
				"00010110" when "00111001", 
				"01010000" when "00111010", 
				"10110101" when "00111011", 
				"11011100" when "00111100", 
				"00111001" when "00111101", 
				"01111111" when "00111110", 
				"10011010" when "00111111", 
				"00100010" when "01000000", 
				"11000111" when "01000001", 
				"10000001" when "01000010", 
				"01100100" when "01000011", 
				"00001101" when "01000100", 
				"11101000" when "01000101", 
				"10101110" when "01000110", 
				"01001011" when "01000111", 
				"01111100" when "01001000", 
				"10011001" when "01001001", 
				"11011111" when "01001010", 
				"00111010" when "01001011", 
				"01010011" when "01001100", 
				"10110110" when "01001101", 
				"11110000" when "01001110", 
				"00010101" when "01001111", 
				"10011110" when "01010000", 
				"01111011" when "01010001", 
				"00111101" when "01010010", 
				"11011000" when "01010011", 
				"10110001" when "01010100", 
				"01010100" when "01010101", 
				"00010010" when "01010110", 
				"11110111" when "01010111", 
				"11000000" when "01011000", 
				"00100101" when "01011001", 
				"01100011" when "01011010", 
				"10000110" when "01011011", 
				"11101111" when "01011100", 
				"00001010" when "01011101", 
				"01001100" when "01011110", 
				"10101001" when "01011111", 
				"00110011" when "01100000", 
				"11010110" when "01100001", 
				"10010000" when "01100010", 
				"01110101" when "01100011", 
				"00011100" when "01100100", 
				"11111001" when "01100101", 
				"10111111" when "01100110", 
				"01011010" when "01100111", 
				"01101101" when "01101000", 
				"10001000" when "01101001", 
				"11001110" when "01101010", 
				"00101011" when "01101011", 
				"01000010" when "01101100", 
				"10100111" when "01101101", 
				"11100001" when "01101110", 
				"00000100" when "01101111", 
				"10001111" when "01110000", 
				"01101010" when "01110001", 
				"00101100" when "01110010", 
				"11001001" when "01110011", 
				"10100000" when "01110100", 
				"01000101" when "01110101", 
				"00000011" when "01110110", 
				"11100110" when "01110111", 
				"11010001" when "01111000", 
				"00110100" when "01111001", 
				"01110010" when "01111010", 
				"10010111" when "01111011", 
				"11111110" when "01111100", 
				"00011011" when "01111101", 
				"01011101" when "01111110", 
				"10111000" when "01111111", 
				"01000100" when "10000000", 
				"10100001" when "10000001", 
				"11100111" when "10000010", 
				"00000010" when "10000011", 
				"01101011" when "10000100", 
				"10001110" when "10000101", 
				"11001000" when "10000110", 
				"00101101" when "10000111", 
				"00011010" when "10001000", 
				"11111111" when "10001001", 
				"10111001" when "10001010", 
				"01011100" when "10001011", 
				"00110101" when "10001100", 
				"11010000" when "10001101", 
				"10010110" when "10001110", 
				"01110011" when "10001111", 
				"11111000" when "10010000", 
				"00011101" when "10010001", 
				"01011011" when "10010010", 
				"10111110" when "10010011", 
				"11010111" when "10010100", 
				"00110010" when "10010101", 
				"01110100" when "10010110", 
				"10010001" when "10010111", 
				"10100110" when "10011000", 
				"01000011" when "10011001", 
				"00000101" when "10011010", 
				"11100000" when "10011011", 
				"10001001" when "10011100", 
				"01101100" when "10011101", 
				"00101010" when "10011110", 
				"11001111" when "10011111", 
				"01010101" when "10100000", 
				"10110000" when "10100001", 
				"11110110" when "10100010", 
				"00010011" when "10100011", 
				"01111010" when "10100100", 
				"10011111" when "10100101", 
				"11011001" when "10100110", 
				"00111100" when "10100111", 
				"00001011" when "10101000", 
				"11101110" when "10101001", 
				"10101000" when "10101010", 
				"01001101" when "10101011", 
				"00100100" when "10101100", 
				"11000001" when "10101101", 
				"10000111" when "10101110", 
				"01100010" when "10101111", 
				"11101001" when "10110000", 
				"00001100" when "10110001", 
				"01001010" when "10110010", 
				"10101111" when "10110011", 
				"11000110" when "10110100", 
				"00100011" when "10110101", 
				"01100101" when "10110110", 
				"10000000" when "10110111", 
				"10110111" when "10111000", 
				"01010010" when "10111001", 
				"00010100" when "10111010", 
				"11110001" when "10111011", 
				"10011000" when "10111100", 
				"01111101" when "10111101", 
				"00111011" when "10111110", 
				"11011110" when "10111111", 
				"01100110" when "11000000", 
				"10000011" when "11000001", 
				"11000101" when "11000010", 
				"00100000" when "11000011", 
				"01001001" when "11000100", 
				"10101100" when "11000101", 
				"11101010" when "11000110", 
				"00001111" when "11000111", 
				"00111000" when "11001000", 
				"11011101" when "11001001", 
				"10011011" when "11001010", 
				"01111110" when "11001011", 
				"00010111" when "11001100", 
				"11110010" when "11001101", 
				"10110100" when "11001110", 
				"01010001" when "11001111", 
				"11011010" when "11010000", 
				"00111111" when "11010001", 
				"01111001" when "11010010", 
				"10011100" when "11010011", 
				"11110101" when "11010100", 
				"00010000" when "11010101", 
				"01010110" when "11010110", 
				"10110011" when "11010111", 
				"10000100" when "11011000", 
				"01100001" when "11011001", 
				"00100111" when "11011010", 
				"11000010" when "11011011", 
				"10101011" when "11011100", 
				"01001110" when "11011101", 
				"00001000" when "11011110", 
				"11101101" when "11011111", 
				"01110111" when "11100000", 
				"10010010" when "11100001", 
				"11010100" when "11100010", 
				"00110001" when "11100011", 
				"01011000" when "11100100", 
				"10111101" when "11100101", 
				"11111011" when "11100110", 
				"00011110" when "11100111", 
				"00101001" when "11101000", 
				"11001100" when "11101001", 
				"10001010" when "11101010", 
				"01101111" when "11101011", 
				"00000110" when "11101100", 
				"11100011" when "11101101", 
				"10100101" when "11101110", 
				"01000000" when "11101111", 
				"11001011" when "11110000", 
				"00101110" when "11110001", 
				"01101000" when "11110010", 
				"10001101" when "11110011", 
				"11100100" when "11110100", 
				"00000001" when "11110101", 
				"01000111" when "11110110", 
				"10100010" when "11110111", 
				"10010101" when "11111000", 
				"01110000" when "11111001", 
				"00110110" when "11111010", 
				"11010011" when "11111011", 
				"10111010" when "11111100", 
				"01011111" when "11111101", 
				"00011001" when "11111110", 
				"11111100" when "11111111";

end mul_E5_mem;

