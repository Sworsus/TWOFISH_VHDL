----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:25:29 04/23/2021 
-- Design Name: 
-- Module Name:    mul_3D_mem - mul_3D_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_3D_mem is
	port (
			in_3D : in STD_LOGIC_VECTOR (7 downto 0);
			out_3D : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_3D_mem;

architecture mul_3D_mem of mul_3D_mem is

begin

	with in_3D select
		out_3D <= "00000000" when "00000000", 
					"00111101" when "00000001", 
					"01111010" when "00000010", 
					"01000111" when "00000011", 
					"11110100" when "00000100", 
					"11001001" when "00000101", 
					"10001110" when "00000110", 
					"10110011" when "00000111", 
					"10000001" when "00001000", 
					"10111100" when "00001001", 
					"11111011" when "00001010", 
					"11000110" when "00001011", 
					"01110101" when "00001100", 
					"01001000" when "00001101", 
					"00001111" when "00001110", 
					"00110010" when "00001111", 
					"01101011" when "00010000", 
					"01010110" when "00010001", 
					"00010001" when "00010010", 
					"00101100" when "00010011", 
					"10011111" when "00010100", 
					"10100010" when "00010101", 
					"11100101" when "00010110", 
					"11011000" when "00010111", 
					"11101010" when "00011000", 
					"11010111" when "00011001", 
					"10010000" when "00011010", 
					"10101101" when "00011011", 
					"00011110" when "00011100", 
					"00100011" when "00011101", 
					"01100100" when "00011110", 
					"01011001" when "00011111", 
					"11010110" when "00100000", 
					"11101011" when "00100001", 
					"10101100" when "00100010", 
					"10010001" when "00100011", 
					"00100010" when "00100100", 
					"00011111" when "00100101", 
					"01011000" when "00100110", 
					"01100101" when "00100111", 
					"01010111" when "00101000", 
					"01101010" when "00101001", 
					"00101101" when "00101010", 
					"00010000" when "00101011", 
					"10100011" when "00101100", 
					"10011110" when "00101101", 
					"11011001" when "00101110", 
					"11100100" when "00101111", 
					"10111101" when "00110000", 
					"10000000" when "00110001", 
					"11000111" when "00110010", 
					"11111010" when "00110011", 
					"01001001" when "00110100", 
					"01110100" when "00110101", 
					"00110011" when "00110110", 
					"00001110" when "00110111", 
					"00111100" when "00111000", 
					"00000001" when "00111001", 
					"01000110" when "00111010", 
					"01111011" when "00111011", 
					"11001000" when "00111100", 
					"11110101" when "00111101", 
					"10110010" when "00111110", 
					"10001111" when "00111111", 
					"11000101" when "01000000", 
					"11111000" when "01000001", 
					"10111111" when "01000010", 
					"10000010" when "01000011", 
					"00110001" when "01000100", 
					"00001100" when "01000101", 
					"01001011" when "01000110", 
					"01110110" when "01000111", 
					"01000100" when "01001000", 
					"01111001" when "01001001", 
					"00111110" when "01001010", 
					"00000011" when "01001011", 
					"10110000" when "01001100", 
					"10001101" when "01001101", 
					"11001010" when "01001110", 
					"11110111" when "01001111", 
					"10101110" when "01010000", 
					"10010011" when "01010001", 
					"11010100" when "01010010", 
					"11101001" when "01010011", 
					"01011010" when "01010100", 
					"01100111" when "01010101", 
					"00100000" when "01010110", 
					"00011101" when "01010111", 
					"00101111" when "01011000", 
					"00010010" when "01011001", 
					"01010101" when "01011010", 
					"01101000" when "01011011", 
					"11011011" when "01011100", 
					"11100110" when "01011101", 
					"10100001" when "01011110", 
					"10011100" when "01011111", 
					"00010011" when "01100000", 
					"00101110" when "01100001", 
					"01101001" when "01100010", 
					"01010100" when "01100011", 
					"11100111" when "01100100", 
					"11011010" when "01100101", 
					"10011101" when "01100110", 
					"10100000" when "01100111", 
					"10010010" when "01101000", 
					"10101111" when "01101001", 
					"11101000" when "01101010", 
					"11010101" when "01101011", 
					"01100110" when "01101100", 
					"01011011" when "01101101", 
					"00011100" when "01101110", 
					"00100001" when "01101111", 
					"01111000" when "01110000", 
					"01000101" when "01110001", 
					"00000010" when "01110010", 
					"00111111" when "01110011", 
					"10001100" when "01110100", 
					"10110001" when "01110101", 
					"11110110" when "01110110", 
					"11001011" when "01110111", 
					"11111001" when "01111000", 
					"11000100" when "01111001", 
					"10000011" when "01111010", 
					"10111110" when "01111011", 
					"00001101" when "01111100", 
					"00110000" when "01111101", 
					"01110111" when "01111110", 
					"01001010" when "01111111", 
					"11100011" when "10000000", 
					"11011110" when "10000001", 
					"10011001" when "10000010", 
					"10100100" when "10000011", 
					"00010111" when "10000100", 
					"00101010" when "10000101", 
					"01101101" when "10000110", 
					"01010000" when "10000111", 
					"01100010" when "10001000", 
					"01011111" when "10001001", 
					"00011000" when "10001010", 
					"00100101" when "10001011", 
					"10010110" when "10001100", 
					"10101011" when "10001101", 
					"11101100" when "10001110", 
					"11010001" when "10001111", 
					"10001000" when "10010000", 
					"10110101" when "10010001", 
					"11110010" when "10010010", 
					"11001111" when "10010011", 
					"01111100" when "10010100", 
					"01000001" when "10010101", 
					"00000110" when "10010110", 
					"00111011" when "10010111", 
					"00001001" when "10011000", 
					"00110100" when "10011001", 
					"01110011" when "10011010", 
					"01001110" when "10011011", 
					"11111101" when "10011100", 
					"11000000" when "10011101", 
					"10000111" when "10011110", 
					"10111010" when "10011111", 
					"00110101" when "10100000", 
					"00001000" when "10100001", 
					"01001111" when "10100010", 
					"01110010" when "10100011", 
					"11000001" when "10100100", 
					"11111100" when "10100101", 
					"10111011" when "10100110", 
					"10000110" when "10100111", 
					"10110100" when "10101000", 
					"10001001" when "10101001", 
					"11001110" when "10101010", 
					"11110011" when "10101011", 
					"01000000" when "10101100", 
					"01111101" when "10101101", 
					"00111010" when "10101110", 
					"00000111" when "10101111", 
					"01011110" when "10110000", 
					"01100011" when "10110001", 
					"00100100" when "10110010", 
					"00011001" when "10110011", 
					"10101010" when "10110100", 
					"10010111" when "10110101", 
					"11010000" when "10110110", 
					"11101101" when "10110111", 
					"11011111" when "10111000", 
					"11100010" when "10111001", 
					"10100101" when "10111010", 
					"10011000" when "10111011", 
					"00101011" when "10111100", 
					"00010110" when "10111101", 
					"01010001" when "10111110", 
					"01101100" when "10111111", 
					"00100110" when "11000000", 
					"00011011" when "11000001", 
					"01011100" when "11000010", 
					"01100001" when "11000011", 
					"11010010" when "11000100", 
					"11101111" when "11000101", 
					"10101000" when "11000110", 
					"10010101" when "11000111", 
					"10100111" when "11001000", 
					"10011010" when "11001001", 
					"11011101" when "11001010", 
					"11100000" when "11001011", 
					"01010011" when "11001100", 
					"01101110" when "11001101", 
					"00101001" when "11001110", 
					"00010100" when "11001111", 
					"01001101" when "11010000", 
					"01110000" when "11010001", 
					"00110111" when "11010010", 
					"00001010" when "11010011", 
					"10111001" when "11010100", 
					"10000100" when "11010101", 
					"11000011" when "11010110", 
					"11111110" when "11010111", 
					"11001100" when "11011000", 
					"11110001" when "11011001", 
					"10110110" when "11011010", 
					"10001011" when "11011011", 
					"00111000" when "11011100", 
					"00000101" when "11011101", 
					"01000010" when "11011110", 
					"01111111" when "11011111", 
					"11110000" when "11100000", 
					"11001101" when "11100001", 
					"10001010" when "11100010", 
					"10110111" when "11100011", 
					"00000100" when "11100100", 
					"00111001" when "11100101", 
					"01111110" when "11100110", 
					"01000011" when "11100111", 
					"01110001" when "11101000", 
					"01001100" when "11101001", 
					"00001011" when "11101010", 
					"00110110" when "11101011", 
					"10000101" when "11101100", 
					"10111000" when "11101101", 
					"11111111" when "11101110", 
					"11000010" when "11101111", 
					"10011011" when "11110000", 
					"10100110" when "11110001", 
					"11100001" when "11110010", 
					"11011100" when "11110011", 
					"01101111" when "11110100", 
					"01010010" when "11110101", 
					"00010101" when "11110110", 
					"00101000" when "11110111", 
					"00011010" when "11111000", 
					"00100111" when "11111001", 
					"01100000" when "11111010", 
					"01011101" when "11111011", 
					"11101110" when "11111100", 
					"11010011" when "11111101", 
					"10010100" when "11111110", 
					"10101001" when "11111111";

end mul_3D_mem;

