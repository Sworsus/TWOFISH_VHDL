----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:14:08 04/24/2021 
-- Design Name: 
-- Module Name:    mul_FC_mem - mul_FC_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_FC_mem is
	port (
			in_FC : in STD_LOGIC_VECTOR (7 downto 0);
			out_FC : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_FC_mem;

architecture mul_FC_mem of mul_FC_mem is

begin

	with in_FC select
	out_FC <= "00000000" when "00000000", 
				"11111100" when "00000001", 
				"10010001" when "00000010", 
				"01101101" when "00000011", 
				"01001011" when "00000100", 
				"10110111" when "00000101", 
				"11011010" when "00000110", 
				"00100110" when "00000111", 
				"10010110" when "00001000", 
				"01101010" when "00001001", 
				"00000111" when "00001010", 
				"11111011" when "00001011", 
				"11011101" when "00001100", 
				"00100001" when "00001101", 
				"01001100" when "00001110", 
				"10110000" when "00001111", 
				"01000101" when "00010000", 
				"10111001" when "00010001", 
				"11010100" when "00010010", 
				"00101000" when "00010011", 
				"00001110" when "00010100", 
				"11110010" when "00010101", 
				"10011111" when "00010110", 
				"01100011" when "00010111", 
				"11010011" when "00011000", 
				"00101111" when "00011001", 
				"01000010" when "00011010", 
				"10111110" when "00011011", 
				"10011000" when "00011100", 
				"01100100" when "00011101", 
				"00001001" when "00011110", 
				"11110101" when "00011111", 
				"10001010" when "00100000", 
				"01110110" when "00100001", 
				"00011011" when "00100010", 
				"11100111" when "00100011", 
				"11000001" when "00100100", 
				"00111101" when "00100101", 
				"01010000" when "00100110", 
				"10101100" when "00100111", 
				"00011100" when "00101000", 
				"11100000" when "00101001", 
				"10001101" when "00101010", 
				"01110001" when "00101011", 
				"01010111" when "00101100", 
				"10101011" when "00101101", 
				"11000110" when "00101110", 
				"00111010" when "00101111", 
				"11001111" when "00110000", 
				"00110011" when "00110001", 
				"01011110" when "00110010", 
				"10100010" when "00110011", 
				"10000100" when "00110100", 
				"01111000" when "00110101", 
				"00010101" when "00110110", 
				"11101001" when "00110111", 
				"01011001" when "00111000", 
				"10100101" when "00111001", 
				"11001000" when "00111010", 
				"00110100" when "00111011", 
				"00010010" when "00111100", 
				"11101110" when "00111101", 
				"10000011" when "00111110", 
				"01111111" when "00111111", 
				"01111101" when "01000000", 
				"10000001" when "01000001", 
				"11101100" when "01000010", 
				"00010000" when "01000011", 
				"00110110" when "01000100", 
				"11001010" when "01000101", 
				"10100111" when "01000110", 
				"01011011" when "01000111", 
				"11101011" when "01001000", 
				"00010111" when "01001001", 
				"01111010" when "01001010", 
				"10000110" when "01001011", 
				"10100000" when "01001100", 
				"01011100" when "01001101", 
				"00110001" when "01001110", 
				"11001101" when "01001111", 
				"00111000" when "01010000", 
				"11000100" when "01010001", 
				"10101001" when "01010010", 
				"01010101" when "01010011", 
				"01110011" when "01010100", 
				"10001111" when "01010101", 
				"11100010" when "01010110", 
				"00011110" when "01010111", 
				"10101110" when "01011000", 
				"01010010" when "01011001", 
				"00111111" when "01011010", 
				"11000011" when "01011011", 
				"11100101" when "01011100", 
				"00011001" when "01011101", 
				"01110100" when "01011110", 
				"10001000" when "01011111", 
				"11110111" when "01100000", 
				"00001011" when "01100001", 
				"01100110" when "01100010", 
				"10011010" when "01100011", 
				"10111100" when "01100100", 
				"01000000" when "01100101", 
				"00101101" when "01100110", 
				"11010001" when "01100111", 
				"01100001" when "01101000", 
				"10011101" when "01101001", 
				"11110000" when "01101010", 
				"00001100" when "01101011", 
				"00101010" when "01101100", 
				"11010110" when "01101101", 
				"10111011" when "01101110", 
				"01000111" when "01101111", 
				"10110010" when "01110000", 
				"01001110" when "01110001", 
				"00100011" when "01110010", 
				"11011111" when "01110011", 
				"11111001" when "01110100", 
				"00000101" when "01110101", 
				"01101000" when "01110110", 
				"10010100" when "01110111", 
				"00100100" when "01111000", 
				"11011000" when "01111001", 
				"10110101" when "01111010", 
				"01001001" when "01111011", 
				"01101111" when "01111100", 
				"10010011" when "01111101", 
				"11111110" when "01111110", 
				"00000010" when "01111111", 
				"11111010" when "10000000", 
				"00000110" when "10000001", 
				"01101011" when "10000010", 
				"10010111" when "10000011", 
				"10110001" when "10000100", 
				"01001101" when "10000101", 
				"00100000" when "10000110", 
				"11011100" when "10000111", 
				"01101100" when "10001000", 
				"10010000" when "10001001", 
				"11111101" when "10001010", 
				"00000001" when "10001011", 
				"00100111" when "10001100", 
				"11011011" when "10001101", 
				"10110110" when "10001110", 
				"01001010" when "10001111", 
				"10111111" when "10010000", 
				"01000011" when "10010001", 
				"00101110" when "10010010", 
				"11010010" when "10010011", 
				"11110100" when "10010100", 
				"00001000" when "10010101", 
				"01100101" when "10010110", 
				"10011001" when "10010111", 
				"00101001" when "10011000", 
				"11010101" when "10011001", 
				"10111000" when "10011010", 
				"01000100" when "10011011", 
				"01100010" when "10011100", 
				"10011110" when "10011101", 
				"11110011" when "10011110", 
				"00001111" when "10011111", 
				"01110000" when "10100000", 
				"10001100" when "10100001", 
				"11100001" when "10100010", 
				"00011101" when "10100011", 
				"00111011" when "10100100", 
				"11000111" when "10100101", 
				"10101010" when "10100110", 
				"01010110" when "10100111", 
				"11100110" when "10101000", 
				"00011010" when "10101001", 
				"01110111" when "10101010", 
				"10001011" when "10101011", 
				"10101101" when "10101100", 
				"01010001" when "10101101", 
				"00111100" when "10101110", 
				"11000000" when "10101111", 
				"00110101" when "10110000", 
				"11001001" when "10110001", 
				"10100100" when "10110010", 
				"01011000" when "10110011", 
				"01111110" when "10110100", 
				"10000010" when "10110101", 
				"11101111" when "10110110", 
				"00010011" when "10110111", 
				"10100011" when "10111000", 
				"01011111" when "10111001", 
				"00110010" when "10111010", 
				"11001110" when "10111011", 
				"11101000" when "10111100", 
				"00010100" when "10111101", 
				"01111001" when "10111110", 
				"10000101" when "10111111", 
				"10000111" when "11000000", 
				"01111011" when "11000001", 
				"00010110" when "11000010", 
				"11101010" when "11000011", 
				"11001100" when "11000100", 
				"00110000" when "11000101", 
				"01011101" when "11000110", 
				"10100001" when "11000111", 
				"00010001" when "11001000", 
				"11101101" when "11001001", 
				"10000000" when "11001010", 
				"01111100" when "11001011", 
				"01011010" when "11001100", 
				"10100110" when "11001101", 
				"11001011" when "11001110", 
				"00110111" when "11001111", 
				"11000010" when "11010000", 
				"00111110" when "11010001", 
				"01010011" when "11010010", 
				"10101111" when "11010011", 
				"10001001" when "11010100", 
				"01110101" when "11010101", 
				"00011000" when "11010110", 
				"11100100" when "11010111", 
				"01010100" when "11011000", 
				"10101000" when "11011001", 
				"11000101" when "11011010", 
				"00111001" when "11011011", 
				"00011111" when "11011100", 
				"11100011" when "11011101", 
				"10001110" when "11011110", 
				"01110010" when "11011111", 
				"00001101" when "11100000", 
				"11110001" when "11100001", 
				"10011100" when "11100010", 
				"01100000" when "11100011", 
				"01000110" when "11100100", 
				"10111010" when "11100101", 
				"11010111" when "11100110", 
				"00101011" when "11100111", 
				"10011011" when "11101000", 
				"01100111" when "11101001", 
				"00001010" when "11101010", 
				"11110110" when "11101011", 
				"11010000" when "11101100", 
				"00101100" when "11101101", 
				"01000001" when "11101110", 
				"10111101" when "11101111", 
				"01001000" when "11110000", 
				"10110100" when "11110001", 
				"11011001" when "11110010", 
				"00100101" when "11110011", 
				"00000011" when "11110100", 
				"11111111" when "11110101", 
				"10010010" when "11110110", 
				"01101110" when "11110111", 
				"11011110" when "11111000", 
				"00100010" when "11111001", 
				"01001111" when "11111010", 
				"10110011" when "11111011", 
				"10010101" when "11111100", 
				"01101001" when "11111101", 
				"00000100" when "11111110", 
				"11111000" when "11111111";

end mul_FC_mem;

