----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:45:57 04/24/2021 
-- Design Name: 
-- Module Name:    mul_9E_mem - mul_9E_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_9E_mem is
	port (
			in_9E : in STD_LOGIC_VECTOR (7 downto 0);
			out_9E : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_9E_mem;

architecture mul_9E_mem of mul_9E_mem is

begin

	with in_9E select
	out_9E <= "00000000" when "00000000", 
				"10011110" when "00000001", 
				"01010101" when "00000010", 
				"11001011" when "00000011", 
				"10101010" when "00000100", 
				"00110100" when "00000101", 
				"11111111" when "00000110", 
				"01100001" when "00000111", 
				"00111101" when "00001000", 
				"10100011" when "00001001", 
				"01101000" when "00001010", 
				"11110110" when "00001011", 
				"10010111" when "00001100", 
				"00001001" when "00001101", 
				"11000010" when "00001110", 
				"01011100" when "00001111", 
				"01111010" when "00010000", 
				"11100100" when "00010001", 
				"00101111" when "00010010", 
				"10110001" when "00010011", 
				"11010000" when "00010100", 
				"01001110" when "00010101", 
				"10000101" when "00010110", 
				"00011011" when "00010111", 
				"01000111" when "00011000", 
				"11011001" when "00011001", 
				"00010010" when "00011010", 
				"10001100" when "00011011", 
				"11101101" when "00011100", 
				"01110011" when "00011101", 
				"10111000" when "00011110", 
				"00100110" when "00011111", 
				"11110100" when "00100000", 
				"01101010" when "00100001", 
				"10100001" when "00100010", 
				"00111111" when "00100011", 
				"01011110" when "00100100", 
				"11000000" when "00100101", 
				"00001011" when "00100110", 
				"10010101" when "00100111", 
				"11001001" when "00101000", 
				"01010111" when "00101001", 
				"10011100" when "00101010", 
				"00000010" when "00101011", 
				"01100011" when "00101100", 
				"11111101" when "00101101", 
				"00110110" when "00101110", 
				"10101000" when "00101111", 
				"10001110" when "00110000", 
				"00010000" when "00110001", 
				"11011011" when "00110010", 
				"01000101" when "00110011", 
				"00100100" when "00110100", 
				"10111010" when "00110101", 
				"01110001" when "00110110", 
				"11101111" when "00110111", 
				"10110011" when "00111000", 
				"00101101" when "00111001", 
				"11100110" when "00111010", 
				"01111000" when "00111011", 
				"00011001" when "00111100", 
				"10000111" when "00111101", 
				"01001100" when "00111110", 
				"11010010" when "00111111", 
				"10000001" when "01000000", 
				"00011111" when "01000001", 
				"11010100" when "01000010", 
				"01001010" when "01000011", 
				"00101011" when "01000100", 
				"10110101" when "01000101", 
				"01111110" when "01000110", 
				"11100000" when "01000111", 
				"10111100" when "01001000", 
				"00100010" when "01001001", 
				"11101001" when "01001010", 
				"01110111" when "01001011", 
				"00010110" when "01001100", 
				"10001000" when "01001101", 
				"01000011" when "01001110", 
				"11011101" when "01001111", 
				"11111011" when "01010000", 
				"01100101" when "01010001", 
				"10101110" when "01010010", 
				"00110000" when "01010011", 
				"01010001" when "01010100", 
				"11001111" when "01010101", 
				"00000100" when "01010110", 
				"10011010" when "01010111", 
				"11000110" when "01011000", 
				"01011000" when "01011001", 
				"10010011" when "01011010", 
				"00001101" when "01011011", 
				"01101100" when "01011100", 
				"11110010" when "01011101", 
				"00111001" when "01011110", 
				"10100111" when "01011111", 
				"01110101" when "01100000", 
				"11101011" when "01100001", 
				"00100000" when "01100010", 
				"10111110" when "01100011", 
				"11011111" when "01100100", 
				"01000001" when "01100101", 
				"10001010" when "01100110", 
				"00010100" when "01100111", 
				"01001000" when "01101000", 
				"11010110" when "01101001", 
				"00011101" when "01101010", 
				"10000011" when "01101011", 
				"11100010" when "01101100", 
				"01111100" when "01101101", 
				"10110111" when "01101110", 
				"00101001" when "01101111", 
				"00001111" when "01110000", 
				"10010001" when "01110001", 
				"01011010" when "01110010", 
				"11000100" when "01110011", 
				"10100101" when "01110100", 
				"00111011" when "01110101", 
				"11110000" when "01110110", 
				"01101110" when "01110111", 
				"00110010" when "01111000", 
				"10101100" when "01111001", 
				"01100111" when "01111010", 
				"11111001" when "01111011", 
				"10011000" when "01111100", 
				"00000110" when "01111101", 
				"11001101" when "01111110", 
				"01010011" when "01111111", 
				"01101011" when "10000000", 
				"11110101" when "10000001", 
				"00111110" when "10000010", 
				"10100000" when "10000011", 
				"11000001" when "10000100", 
				"01011111" when "10000101", 
				"10010100" when "10000110", 
				"00001010" when "10000111", 
				"01010110" when "10001000", 
				"11001000" when "10001001", 
				"00000011" when "10001010", 
				"10011101" when "10001011", 
				"11111100" when "10001100", 
				"01100010" when "10001101", 
				"10101001" when "10001110", 
				"00110111" when "10001111", 
				"00010001" when "10010000", 
				"10001111" when "10010001", 
				"01000100" when "10010010", 
				"11011010" when "10010011", 
				"10111011" when "10010100", 
				"00100101" when "10010101", 
				"11101110" when "10010110", 
				"01110000" when "10010111", 
				"00101100" when "10011000", 
				"10110010" when "10011001", 
				"01111001" when "10011010", 
				"11100111" when "10011011", 
				"10000110" when "10011100", 
				"00011000" when "10011101", 
				"11010011" when "10011110", 
				"01001101" when "10011111", 
				"10011111" when "10100000", 
				"00000001" when "10100001", 
				"11001010" when "10100010", 
				"01010100" when "10100011", 
				"00110101" when "10100100", 
				"10101011" when "10100101", 
				"01100000" when "10100110", 
				"11111110" when "10100111", 
				"10100010" when "10101000", 
				"00111100" when "10101001", 
				"11110111" when "10101010", 
				"01101001" when "10101011", 
				"00001000" when "10101100", 
				"10010110" when "10101101", 
				"01011101" when "10101110", 
				"11000011" when "10101111", 
				"11100101" when "10110000", 
				"01111011" when "10110001", 
				"10110000" when "10110010", 
				"00101110" when "10110011", 
				"01001111" when "10110100", 
				"11010001" when "10110101", 
				"00011010" when "10110110", 
				"10000100" when "10110111", 
				"11011000" when "10111000", 
				"01000110" when "10111001", 
				"10001101" when "10111010", 
				"00010011" when "10111011", 
				"01110010" when "10111100", 
				"11101100" when "10111101", 
				"00100111" when "10111110", 
				"10111001" when "10111111", 
				"11101010" when "11000000", 
				"01110100" when "11000001", 
				"10111111" when "11000010", 
				"00100001" when "11000011", 
				"01000000" when "11000100", 
				"11011110" when "11000101", 
				"00010101" when "11000110", 
				"10001011" when "11000111", 
				"11010111" when "11001000", 
				"01001001" when "11001001", 
				"10000010" when "11001010", 
				"00011100" when "11001011", 
				"01111101" when "11001100", 
				"11100011" when "11001101", 
				"00101000" when "11001110", 
				"10110110" when "11001111", 
				"10010000" when "11010000", 
				"00001110" when "11010001", 
				"11000101" when "11010010", 
				"01011011" when "11010011", 
				"00111010" when "11010100", 
				"10100100" when "11010101", 
				"01101111" when "11010110", 
				"11110001" when "11010111", 
				"10101101" when "11011000", 
				"00110011" when "11011001", 
				"11111000" when "11011010", 
				"01100110" when "11011011", 
				"00000111" when "11011100", 
				"10011001" when "11011101", 
				"01010010" when "11011110", 
				"11001100" when "11011111", 
				"00011110" when "11100000", 
				"10000000" when "11100001", 
				"01001011" when "11100010", 
				"11010101" when "11100011", 
				"10110100" when "11100100", 
				"00101010" when "11100101", 
				"11100001" when "11100110", 
				"01111111" when "11100111", 
				"00100011" when "11101000", 
				"10111101" when "11101001", 
				"01110110" when "11101010", 
				"11101000" when "11101011", 
				"10001001" when "11101100", 
				"00010111" when "11101101", 
				"11011100" when "11101110", 
				"01000010" when "11101111", 
				"01100100" when "11110000", 
				"11111010" when "11110001", 
				"00110001" when "11110010", 
				"10101111" when "11110011", 
				"11001110" when "11110100", 
				"01010000" when "11110101", 
				"10011011" when "11110110", 
				"00000101" when "11110111", 
				"01011001" when "11111000", 
				"11000111" when "11111001", 
				"00001100" when "11111010", 
				"10010010" when "11111011", 
				"11110011" when "11111100", 
				"01101101" when "11111101", 
				"10100110" when "11111110", 
				"00111000" when "11111111";

end mul_9E_mem;

