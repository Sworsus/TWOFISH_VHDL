----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:10:40 04/24/2021 
-- Design Name: 
-- Module Name:    mul_68_mem - mul_68_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_68_mem is
	port (
			in_68 : in STD_LOGIC_VECTOR (7 downto 0);
			out_68 : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_68_mem;

architecture mul_68_mem of mul_68_mem is

begin

	with in_68 select
	out_68 <= "00000000" when "00000000", 
				"01101000" when "00000001", 
				"11010000" when "00000010", 
				"10111000" when "00000011", 
				"11001001" when "00000100", 
				"10100001" when "00000101", 
				"00011001" when "00000110", 
				"01110001" when "00000111", 
				"11111011" when "00001000", 
				"10010011" when "00001001", 
				"00101011" when "00001010", 
				"01000011" when "00001011", 
				"00110010" when "00001100", 
				"01011010" when "00001101", 
				"11100010" when "00001110", 
				"10001010" when "00001111", 
				"10011111" when "00010000", 
				"11110111" when "00010001", 
				"01001111" when "00010010", 
				"00100111" when "00010011", 
				"01010110" when "00010100", 
				"00111110" when "00010101", 
				"10000110" when "00010110", 
				"11101110" when "00010111", 
				"01100100" when "00011000", 
				"00001100" when "00011001", 
				"10110100" when "00011010", 
				"11011100" when "00011011", 
				"10101101" when "00011100", 
				"11000101" when "00011101", 
				"01111101" when "00011110", 
				"00010101" when "00011111", 
				"01010111" when "00100000", 
				"00111111" when "00100001", 
				"10000111" when "00100010", 
				"11101111" when "00100011", 
				"10011110" when "00100100", 
				"11110110" when "00100101", 
				"01001110" when "00100110", 
				"00100110" when "00100111", 
				"10101100" when "00101000", 
				"11000100" when "00101001", 
				"01111100" when "00101010", 
				"00010100" when "00101011", 
				"01100101" when "00101100", 
				"00001101" when "00101101", 
				"10110101" when "00101110", 
				"11011101" when "00101111", 
				"11001000" when "00110000", 
				"10100000" when "00110001", 
				"00011000" when "00110010", 
				"01110000" when "00110011", 
				"00000001" when "00110100", 
				"01101001" when "00110101", 
				"11010001" when "00110110", 
				"10111001" when "00110111", 
				"00110011" when "00111000", 
				"01011011" when "00111001", 
				"11100011" when "00111010", 
				"10001011" when "00111011", 
				"11111010" when "00111100", 
				"10010010" when "00111101", 
				"00101010" when "00111110", 
				"01000010" when "00111111", 
				"10101110" when "01000000", 
				"11000110" when "01000001", 
				"01111110" when "01000010", 
				"00010110" when "01000011", 
				"01100111" when "01000100", 
				"00001111" when "01000101", 
				"10110111" when "01000110", 
				"11011111" when "01000111", 
				"01010101" when "01001000", 
				"00111101" when "01001001", 
				"10000101" when "01001010", 
				"11101101" when "01001011", 
				"10011100" when "01001100", 
				"11110100" when "01001101", 
				"01001100" when "01001110", 
				"00100100" when "01001111", 
				"00110001" when "01010000", 
				"01011001" when "01010001", 
				"11100001" when "01010010", 
				"10001001" when "01010011", 
				"11111000" when "01010100", 
				"10010000" when "01010101", 
				"00101000" when "01010110", 
				"01000000" when "01010111", 
				"11001010" when "01011000", 
				"10100010" when "01011001", 
				"00011010" when "01011010", 
				"01110010" when "01011011", 
				"00000011" when "01011100", 
				"01101011" when "01011101", 
				"11010011" when "01011110", 
				"10111011" when "01011111", 
				"11111001" when "01100000", 
				"10010001" when "01100001", 
				"00101001" when "01100010", 
				"01000001" when "01100011", 
				"00110000" when "01100100", 
				"01011000" when "01100101", 
				"11100000" when "01100110", 
				"10001000" when "01100111", 
				"00000010" when "01101000", 
				"01101010" when "01101001", 
				"11010010" when "01101010", 
				"10111010" when "01101011", 
				"11001011" when "01101100", 
				"10100011" when "01101101", 
				"00011011" when "01101110", 
				"01110011" when "01101111", 
				"01100110" when "01110000", 
				"00001110" when "01110001", 
				"10110110" when "01110010", 
				"11011110" when "01110011", 
				"10101111" when "01110100", 
				"11000111" when "01110101", 
				"01111111" when "01110110", 
				"00010111" when "01110111", 
				"10011101" when "01111000", 
				"11110101" when "01111001", 
				"01001101" when "01111010", 
				"00100101" when "01111011", 
				"01010100" when "01111100", 
				"00111100" when "01111101", 
				"10000100" when "01111110", 
				"11101100" when "01111111", 
				"00110101" when "10000000", 
				"01011101" when "10000001", 
				"11100101" when "10000010", 
				"10001101" when "10000011", 
				"11111100" when "10000100", 
				"10010100" when "10000101", 
				"00101100" when "10000110", 
				"01000100" when "10000111", 
				"11001110" when "10001000", 
				"10100110" when "10001001", 
				"00011110" when "10001010", 
				"01110110" when "10001011", 
				"00000111" when "10001100", 
				"01101111" when "10001101", 
				"11010111" when "10001110", 
				"10111111" when "10001111", 
				"10101010" when "10010000", 
				"11000010" when "10010001", 
				"01111010" when "10010010", 
				"00010010" when "10010011", 
				"01100011" when "10010100", 
				"00001011" when "10010101", 
				"10110011" when "10010110", 
				"11011011" when "10010111", 
				"01010001" when "10011000", 
				"00111001" when "10011001", 
				"10000001" when "10011010", 
				"11101001" when "10011011", 
				"10011000" when "10011100", 
				"11110000" when "10011101", 
				"01001000" when "10011110", 
				"00100000" when "10011111", 
				"01100010" when "10100000", 
				"00001010" when "10100001", 
				"10110010" when "10100010", 
				"11011010" when "10100011", 
				"10101011" when "10100100", 
				"11000011" when "10100101", 
				"01111011" when "10100110", 
				"00010011" when "10100111", 
				"10011001" when "10101000", 
				"11110001" when "10101001", 
				"01001001" when "10101010", 
				"00100001" when "10101011", 
				"01010000" when "10101100", 
				"00111000" when "10101101", 
				"10000000" when "10101110", 
				"11101000" when "10101111", 
				"11111101" when "10110000", 
				"10010101" when "10110001", 
				"00101101" when "10110010", 
				"01000101" when "10110011", 
				"00110100" when "10110100", 
				"01011100" when "10110101", 
				"11100100" when "10110110", 
				"10001100" when "10110111", 
				"00000110" when "10111000", 
				"01101110" when "10111001", 
				"11010110" when "10111010", 
				"10111110" when "10111011", 
				"11001111" when "10111100", 
				"10100111" when "10111101", 
				"00011111" when "10111110", 
				"01110111" when "10111111", 
				"10011011" when "11000000", 
				"11110011" when "11000001", 
				"01001011" when "11000010", 
				"00100011" when "11000011", 
				"01010010" when "11000100", 
				"00111010" when "11000101", 
				"10000010" when "11000110", 
				"11101010" when "11000111", 
				"01100000" when "11001000", 
				"00001000" when "11001001", 
				"10110000" when "11001010", 
				"11011000" when "11001011", 
				"10101001" when "11001100", 
				"11000001" when "11001101", 
				"01111001" when "11001110", 
				"00010001" when "11001111", 
				"00000100" when "11010000", 
				"01101100" when "11010001", 
				"11010100" when "11010010", 
				"10111100" when "11010011", 
				"11001101" when "11010100", 
				"10100101" when "11010101", 
				"00011101" when "11010110", 
				"01110101" when "11010111", 
				"11111111" when "11011000", 
				"10010111" when "11011001", 
				"00101111" when "11011010", 
				"01000111" when "11011011", 
				"00110110" when "11011100", 
				"01011110" when "11011101", 
				"11100110" when "11011110", 
				"10001110" when "11011111", 
				"11001100" when "11100000", 
				"10100100" when "11100001", 
				"00011100" when "11100010", 
				"01110100" when "11100011", 
				"00000101" when "11100100", 
				"01101101" when "11100101", 
				"11010101" when "11100110", 
				"10111101" when "11100111", 
				"00110111" when "11101000", 
				"01011111" when "11101001", 
				"11100111" when "11101010", 
				"10001111" when "11101011", 
				"11111110" when "11101100", 
				"10010110" when "11101101", 
				"00101110" when "11101110", 
				"01000110" when "11101111", 
				"01010011" when "11110000", 
				"00111011" when "11110001", 
				"10000011" when "11110010", 
				"11101011" when "11110011", 
				"10011010" when "11110100", 
				"11110010" when "11110101", 
				"01001010" when "11110110", 
				"00100010" when "11110111", 
				"10101000" when "11111000", 
				"11000000" when "11111001", 
				"01111000" when "11111010", 
				"00010000" when "11111011", 
				"01100001" when "11111100", 
				"00001001" when "11111101", 
				"10110001" when "11111110", 
				"11011001" when "11111111";

end mul_68_mem;

