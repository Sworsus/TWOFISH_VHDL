----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:09:10 04/24/2021 
-- Design Name: 
-- Module Name:    mul_A1_mem - mul_A1_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_A1_mem is
	port (
			in_A1 : in STD_LOGIC_VECTOR (7 downto 0);
			out_A1 : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_A1_mem;

architecture mul_A1_mem of mul_A1_mem is

begin

	with in_A1 select
	out_A1 <= "00000000" when "00000000", 
				"10100001" when "00000001", 
				"00101011" when "00000010", 
				"10001010" when "00000011", 
				"01010110" when "00000100", 
				"11110111" when "00000101", 
				"01111101" when "00000110", 
				"11011100" when "00000111", 
				"10101100" when "00001000", 
				"00001101" when "00001001", 
				"10000111" when "00001010", 
				"00100110" when "00001011", 
				"11111010" when "00001100", 
				"01011011" when "00001101", 
				"11010001" when "00001110", 
				"01110000" when "00001111", 
				"00110001" when "00010000", 
				"10010000" when "00010001", 
				"00011010" when "00010010", 
				"10111011" when "00010011", 
				"01100111" when "00010100", 
				"11000110" when "00010101", 
				"01001100" when "00010110", 
				"11101101" when "00010111", 
				"10011101" when "00011000", 
				"00111100" when "00011001", 
				"10110110" when "00011010", 
				"00010111" when "00011011", 
				"11001011" when "00011100", 
				"01101010" when "00011101", 
				"11100000" when "00011110", 
				"01000001" when "00011111", 
				"01100010" when "00100000", 
				"11000011" when "00100001", 
				"01001001" when "00100010", 
				"11101000" when "00100011", 
				"00110100" when "00100100", 
				"10010101" when "00100101", 
				"00011111" when "00100110", 
				"10111110" when "00100111", 
				"11001110" when "00101000", 
				"01101111" when "00101001", 
				"11100101" when "00101010", 
				"01000100" when "00101011", 
				"10011000" when "00101100", 
				"00111001" when "00101101", 
				"10110011" when "00101110", 
				"00010010" when "00101111", 
				"01010011" when "00110000", 
				"11110010" when "00110001", 
				"01111000" when "00110010", 
				"11011001" when "00110011", 
				"00000101" when "00110100", 
				"10100100" when "00110101", 
				"00101110" when "00110110", 
				"10001111" when "00110111", 
				"11111111" when "00111000", 
				"01011110" when "00111001", 
				"11010100" when "00111010", 
				"01110101" when "00111011", 
				"10101001" when "00111100", 
				"00001000" when "00111101", 
				"10000010" when "00111110", 
				"00100011" when "00111111", 
				"11000100" when "01000000", 
				"01100101" when "01000001", 
				"11101111" when "01000010", 
				"01001110" when "01000011", 
				"10010010" when "01000100", 
				"00110011" when "01000101", 
				"10111001" when "01000110", 
				"00011000" when "01000111", 
				"01101000" when "01001000", 
				"11001001" when "01001001", 
				"01000011" when "01001010", 
				"11100010" when "01001011", 
				"00111110" when "01001100", 
				"10011111" when "01001101", 
				"00010101" when "01001110", 
				"10110100" when "01001111", 
				"11110101" when "01010000", 
				"01010100" when "01010001", 
				"11011110" when "01010010", 
				"01111111" when "01010011", 
				"10100011" when "01010100", 
				"00000010" when "01010101", 
				"10001000" when "01010110", 
				"00101001" when "01010111", 
				"01011001" when "01011000", 
				"11111000" when "01011001", 
				"01110010" when "01011010", 
				"11010011" when "01011011", 
				"00001111" when "01011100", 
				"10101110" when "01011101", 
				"00100100" when "01011110", 
				"10000101" when "01011111", 
				"10100110" when "01100000", 
				"00000111" when "01100001", 
				"10001101" when "01100010", 
				"00101100" when "01100011", 
				"11110000" when "01100100", 
				"01010001" when "01100101", 
				"11011011" when "01100110", 
				"01111010" when "01100111", 
				"00001010" when "01101000", 
				"10101011" when "01101001", 
				"00100001" when "01101010", 
				"10000000" when "01101011", 
				"01011100" when "01101100", 
				"11111101" when "01101101", 
				"01110111" when "01101110", 
				"11010110" when "01101111", 
				"10010111" when "01110000", 
				"00110110" when "01110001", 
				"10111100" when "01110010", 
				"00011101" when "01110011", 
				"11000001" when "01110100", 
				"01100000" when "01110101", 
				"11101010" when "01110110", 
				"01001011" when "01110111", 
				"00111011" when "01111000", 
				"10011010" when "01111001", 
				"00010000" when "01111010", 
				"10110001" when "01111011", 
				"01101101" when "01111100", 
				"11001100" when "01111101", 
				"01000110" when "01111110", 
				"11100111" when "01111111", 
				"11100001" when "10000000", 
				"01000000" when "10000001", 
				"11001010" when "10000010", 
				"01101011" when "10000011", 
				"10110111" when "10000100", 
				"00010110" when "10000101", 
				"10011100" when "10000110", 
				"00111101" when "10000111", 
				"01001101" when "10001000", 
				"11101100" when "10001001", 
				"01100110" when "10001010", 
				"11000111" when "10001011", 
				"00011011" when "10001100", 
				"10111010" when "10001101", 
				"00110000" when "10001110", 
				"10010001" when "10001111", 
				"11010000" when "10010000", 
				"01110001" when "10010001", 
				"11111011" when "10010010", 
				"01011010" when "10010011", 
				"10000110" when "10010100", 
				"00100111" when "10010101", 
				"10101101" when "10010110", 
				"00001100" when "10010111", 
				"01111100" when "10011000", 
				"11011101" when "10011001", 
				"01010111" when "10011010", 
				"11110110" when "10011011", 
				"00101010" when "10011100", 
				"10001011" when "10011101", 
				"00000001" when "10011110", 
				"10100000" when "10011111", 
				"10000011" when "10100000", 
				"00100010" when "10100001", 
				"10101000" when "10100010", 
				"00001001" when "10100011", 
				"11010101" when "10100100", 
				"01110100" when "10100101", 
				"11111110" when "10100110", 
				"01011111" when "10100111", 
				"00101111" when "10101000", 
				"10001110" when "10101001", 
				"00000100" when "10101010", 
				"10100101" when "10101011", 
				"01111001" when "10101100", 
				"11011000" when "10101101", 
				"01010010" when "10101110", 
				"11110011" when "10101111", 
				"10110010" when "10110000", 
				"00010011" when "10110001", 
				"10011001" when "10110010", 
				"00111000" when "10110011", 
				"11100100" when "10110100", 
				"01000101" when "10110101", 
				"11001111" when "10110110", 
				"01101110" when "10110111", 
				"00011110" when "10111000", 
				"10111111" when "10111001", 
				"00110101" when "10111010", 
				"10010100" when "10111011", 
				"01001000" when "10111100", 
				"11101001" when "10111101", 
				"01100011" when "10111110", 
				"11000010" when "10111111", 
				"00100101" when "11000000", 
				"10000100" when "11000001", 
				"00001110" when "11000010", 
				"10101111" when "11000011", 
				"01110011" when "11000100", 
				"11010010" when "11000101", 
				"01011000" when "11000110", 
				"11111001" when "11000111", 
				"10001001" when "11001000", 
				"00101000" when "11001001", 
				"10100010" when "11001010", 
				"00000011" when "11001011", 
				"11011111" when "11001100", 
				"01111110" when "11001101", 
				"11110100" when "11001110", 
				"01010101" when "11001111", 
				"00010100" when "11010000", 
				"10110101" when "11010001", 
				"00111111" when "11010010", 
				"10011110" when "11010011", 
				"01000010" when "11010100", 
				"11100011" when "11010101", 
				"01101001" when "11010110", 
				"11001000" when "11010111", 
				"10111000" when "11011000", 
				"00011001" when "11011001", 
				"10010011" when "11011010", 
				"00110010" when "11011011", 
				"11101110" when "11011100", 
				"01001111" when "11011101", 
				"11000101" when "11011110", 
				"01100100" when "11011111", 
				"01000111" when "11100000", 
				"11100110" when "11100001", 
				"01101100" when "11100010", 
				"11001101" when "11100011", 
				"00010001" when "11100100", 
				"10110000" when "11100101", 
				"00111010" when "11100110", 
				"10011011" when "11100111", 
				"11101011" when "11101000", 
				"01001010" when "11101001", 
				"11000000" when "11101010", 
				"01100001" when "11101011", 
				"10111101" when "11101100", 
				"00011100" when "11101101", 
				"10010110" when "11101110", 
				"00110111" when "11101111", 
				"01110110" when "11110000", 
				"11010111" when "11110001", 
				"01011101" when "11110010", 
				"11111100" when "11110011", 
				"00100000" when "11110100", 
				"10000001" when "11110101", 
				"00001011" when "11110110", 
				"10101010" when "11110111", 
				"11011010" when "11111000", 
				"01111011" when "11111001", 
				"11110001" when "11111010", 
				"01010000" when "11111011", 
				"10001100" when "11111100", 
				"00101101" when "11111101", 
				"10100111" when "11111110", 
				"00000110" when "11111111";

end mul_A1_mem;

