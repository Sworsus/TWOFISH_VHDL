----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:30:22 04/24/2021 
-- Design Name: 
-- Module Name:    mul_AE_mem - mul_AE_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_AE_mem is
	port (
			in_AE : in STD_LOGIC_VECTOR (7 downto 0);
			out_AE : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_AE_mem;

architecture mul_AE_mem of mul_AE_mem is

begin

	with in_AE select
	out_AE <= "00000000" when "00000000", 
				"10101110" when "00000001", 
				"00110101" when "00000010", 
				"10011011" when "00000011", 
				"01101010" when "00000100", 
				"11000100" when "00000101", 
				"01011111" when "00000110", 
				"11110001" when "00000111", 
				"11010100" when "00001000", 
				"01111010" when "00001001", 
				"11100001" when "00001010", 
				"01001111" when "00001011", 
				"10111110" when "00001100", 
				"00010000" when "00001101", 
				"10001011" when "00001110", 
				"00100101" when "00001111", 
				"11000001" when "00010000", 
				"01101111" when "00010001", 
				"11110100" when "00010010", 
				"01011010" when "00010011", 
				"10101011" when "00010100", 
				"00000101" when "00010101", 
				"10011110" when "00010110", 
				"00110000" when "00010111", 
				"00010101" when "00011000", 
				"10111011" when "00011001", 
				"00100000" when "00011010", 
				"10001110" when "00011011", 
				"01111111" when "00011100", 
				"11010001" when "00011101", 
				"01001010" when "00011110", 
				"11100100" when "00011111", 
				"11101011" when "00100000", 
				"01000101" when "00100001", 
				"11011110" when "00100010", 
				"01110000" when "00100011", 
				"10000001" when "00100100", 
				"00101111" when "00100101", 
				"10110100" when "00100110", 
				"00011010" when "00100111", 
				"00111111" when "00101000", 
				"10010001" when "00101001", 
				"00001010" when "00101010", 
				"10100100" when "00101011", 
				"01010101" when "00101100", 
				"11111011" when "00101101", 
				"01100000" when "00101110", 
				"11001110" when "00101111", 
				"00101010" when "00110000", 
				"10000100" when "00110001", 
				"00011111" when "00110010", 
				"10110001" when "00110011", 
				"01000000" when "00110100", 
				"11101110" when "00110101", 
				"01110101" when "00110110", 
				"11011011" when "00110111", 
				"11111110" when "00111000", 
				"01010000" when "00111001", 
				"11001011" when "00111010", 
				"01100101" when "00111011", 
				"10010100" when "00111100", 
				"00111010" when "00111101", 
				"10100001" when "00111110", 
				"00001111" when "00111111", 
				"10111111" when "01000000", 
				"00010001" when "01000001", 
				"10001010" when "01000010", 
				"00100100" when "01000011", 
				"11010101" when "01000100", 
				"01111011" when "01000101", 
				"11100000" when "01000110", 
				"01001110" when "01000111", 
				"01101011" when "01001000", 
				"11000101" when "01001001", 
				"01011110" when "01001010", 
				"11110000" when "01001011", 
				"00000001" when "01001100", 
				"10101111" when "01001101", 
				"00110100" when "01001110", 
				"10011010" when "01001111", 
				"01111110" when "01010000", 
				"11010000" when "01010001", 
				"01001011" when "01010010", 
				"11100101" when "01010011", 
				"00010100" when "01010100", 
				"10111010" when "01010101", 
				"00100001" when "01010110", 
				"10001111" when "01010111", 
				"10101010" when "01011000", 
				"00000100" when "01011001", 
				"10011111" when "01011010", 
				"00110001" when "01011011", 
				"11000000" when "01011100", 
				"01101110" when "01011101", 
				"11110101" when "01011110", 
				"01011011" when "01011111", 
				"01010100" when "01100000", 
				"11111010" when "01100001", 
				"01100001" when "01100010", 
				"11001111" when "01100011", 
				"00111110" when "01100100", 
				"10010000" when "01100101", 
				"00001011" when "01100110", 
				"10100101" when "01100111", 
				"10000000" when "01101000", 
				"00101110" when "01101001", 
				"10110101" when "01101010", 
				"00011011" when "01101011", 
				"11101010" when "01101100", 
				"01000100" when "01101101", 
				"11011111" when "01101110", 
				"01110001" when "01101111", 
				"10010101" when "01110000", 
				"00111011" when "01110001", 
				"10100000" when "01110010", 
				"00001110" when "01110011", 
				"11111111" when "01110100", 
				"01010001" when "01110101", 
				"11001010" when "01110110", 
				"01100100" when "01110111", 
				"01000001" when "01111000", 
				"11101111" when "01111001", 
				"01110100" when "01111010", 
				"11011010" when "01111011", 
				"00101011" when "01111100", 
				"10000101" when "01111101", 
				"00011110" when "01111110", 
				"10110000" when "01111111", 
				"00010111" when "10000000", 
				"10111001" when "10000001", 
				"00100010" when "10000010", 
				"10001100" when "10000011", 
				"01111101" when "10000100", 
				"11010011" when "10000101", 
				"01001000" when "10000110", 
				"11100110" when "10000111", 
				"11000011" when "10001000", 
				"01101101" when "10001001", 
				"11110110" when "10001010", 
				"01011000" when "10001011", 
				"10101001" when "10001100", 
				"00000111" when "10001101", 
				"10011100" when "10001110", 
				"00110010" when "10001111", 
				"11010110" when "10010000", 
				"01111000" when "10010001", 
				"11100011" when "10010010", 
				"01001101" when "10010011", 
				"10111100" when "10010100", 
				"00010010" when "10010101", 
				"10001001" when "10010110", 
				"00100111" when "10010111", 
				"00000010" when "10011000", 
				"10101100" when "10011001", 
				"00110111" when "10011010", 
				"10011001" when "10011011", 
				"01101000" when "10011100", 
				"11000110" when "10011101", 
				"01011101" when "10011110", 
				"11110011" when "10011111", 
				"11111100" when "10100000", 
				"01010010" when "10100001", 
				"11001001" when "10100010", 
				"01100111" when "10100011", 
				"10010110" when "10100100", 
				"00111000" when "10100101", 
				"10100011" when "10100110", 
				"00001101" when "10100111", 
				"00101000" when "10101000", 
				"10000110" when "10101001", 
				"00011101" when "10101010", 
				"10110011" when "10101011", 
				"01000010" when "10101100", 
				"11101100" when "10101101", 
				"01110111" when "10101110", 
				"11011001" when "10101111", 
				"00111101" when "10110000", 
				"10010011" when "10110001", 
				"00001000" when "10110010", 
				"10100110" when "10110011", 
				"01010111" when "10110100", 
				"11111001" when "10110101", 
				"01100010" when "10110110", 
				"11001100" when "10110111", 
				"11101001" when "10111000", 
				"01000111" when "10111001", 
				"11011100" when "10111010", 
				"01110010" when "10111011", 
				"10000011" when "10111100", 
				"00101101" when "10111101", 
				"10110110" when "10111110", 
				"00011000" when "10111111", 
				"10101000" when "11000000", 
				"00000110" when "11000001", 
				"10011101" when "11000010", 
				"00110011" when "11000011", 
				"11000010" when "11000100", 
				"01101100" when "11000101", 
				"11110111" when "11000110", 
				"01011001" when "11000111", 
				"01111100" when "11001000", 
				"11010010" when "11001001", 
				"01001001" when "11001010", 
				"11100111" when "11001011", 
				"00010110" when "11001100", 
				"10111000" when "11001101", 
				"00100011" when "11001110", 
				"10001101" when "11001111", 
				"01101001" when "11010000", 
				"11000111" when "11010001", 
				"01011100" when "11010010", 
				"11110010" when "11010011", 
				"00000011" when "11010100", 
				"10101101" when "11010101", 
				"00110110" when "11010110", 
				"10011000" when "11010111", 
				"10111101" when "11011000", 
				"00010011" when "11011001", 
				"10001000" when "11011010", 
				"00100110" when "11011011", 
				"11010111" when "11011100", 
				"01111001" when "11011101", 
				"11100010" when "11011110", 
				"01001100" when "11011111", 
				"01000011" when "11100000", 
				"11101101" when "11100001", 
				"01110110" when "11100010", 
				"11011000" when "11100011", 
				"00101001" when "11100100", 
				"10000111" when "11100101", 
				"00011100" when "11100110", 
				"10110010" when "11100111", 
				"10010111" when "11101000", 
				"00111001" when "11101001", 
				"10100010" when "11101010", 
				"00001100" when "11101011", 
				"11111101" when "11101100", 
				"01010011" when "11101101", 
				"11001000" when "11101110", 
				"01100110" when "11101111", 
				"10000010" when "11110000", 
				"00101100" when "11110001", 
				"10110111" when "11110010", 
				"00011001" when "11110011", 
				"11101000" when "11110100", 
				"01000110" when "11110101", 
				"11011101" when "11110110", 
				"01110011" when "11110111", 
				"01010110" when "11111000", 
				"11111000" when "11111001", 
				"01100011" when "11111010", 
				"11001101" when "11111011", 
				"00111100" when "11111100", 
				"10010010" when "11111101", 
				"00001001" when "11111110", 
				"10100111" when "11111111";

end mul_AE_mem;

