----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:52:58 04/23/2021 
-- Design Name: 
-- Module Name:    mul_03_mem - mul_03_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_03_mem is
	port	(
			in_03	: in STD_LOGIC_VECTOR(7 DOWNTO 0);
			out_03 : out STD_LOGIC_VECTOR(7 DOWNTO 0)
			);
end mul_03_mem;

architecture mul_03_mem of mul_03_mem is

begin

	with in_03 select
		out_03 <= "00000000" when "00000000", "00000011" when "00000001", "00000110" when "00000010", "00000101" when "00000011", 
					"00001100" when "00000100", "00001111" when "00000101", "00001010" when "00000110", "00001001" when "00000111", 
					"00011000" when "00001000", "00011011" when "00001001", "00011110" when "00001010", "00011101" when "00001011", 
					"00010100" when "00001100", "00010111" when "00001101", "00010010" when "00001110", "00010001" when "00001111", 
					"00110000" when "00010000", "00110011" when "00010001", "00110110" when "00010010", "00110101" when "00010011", 
					"00111100" when "00010100", "00111111" when "00010101", "00111010" when "00010110", "00111001" when "00010111", 
					"00101000" when "00011000", "00101011" when "00011001", "00101110" when "00011010", "00101101" when "00011011", 
					"00100100" when "00011100", "00100111" when "00011101", "00100010" when "00011110", "00100001" when "00011111", 
					"01100000" when "00100000", "01100011" when "00100001", "01100110" when "00100010", "01100101" when "00100011", 
					"01101100" when "00100100", "01101111" when "00100101", "01101010" when "00100110", "01101001" when "00100111", 
					"01111000" when "00101000", "01111011" when "00101001", "01111110" when "00101010", "01111101" when "00101011", 
					"01110100" when "00101100", "01110111" when "00101101", "01110010" when "00101110", "01110001" when "00101111", 
					"01010000" when "00110000", "01010011" when "00110001", "01010110" when "00110010", "01010101" when "00110011", 
					"01011100" when "00110100", "01011111" when "00110101", "01011010" when "00110110", "01011001" when "00110111", 
					"01001000" when "00111000", "01001011" when "00111001", "01001110" when "00111010", "01001101" when "00111011", 
					"01000100" when "00111100", "01000111" when "00111101", "01000010" when "00111110", "01000001" when "00111111", 
					"11000000" when "01000000", "11000011" when "01000001", "11000110" when "01000010", "11000101" when "01000011", 
					"11001100" when "01000100", "11001111" when "01000101", "11001010" when "01000110", "11001001" when "01000111", 
					"11011000" when "01001000", "11011011" when "01001001", "11011110" when "01001010", "11011101" when "01001011", 
					"11010100" when "01001100", "11010111" when "01001101", "11010010" when "01001110", "11010001" when "01001111", 
					"11110000" when "01010000", "11110011" when "01010001", "11110110" when "01010010", "11110101" when "01010011", 
					"11111100" when "01010100", "11111111" when "01010101", "11111010" when "01010110", "11111001" when "01010111", 
					"11101000" when "01011000", "11101011" when "01011001", "11101110" when "01011010", "11101101" when "01011011", 
					"11100100" when "01011100", "11100111" when "01011101", "11100010" when "01011110", "11100001" when "01011111", 
					"10100000" when "01100000", "10100011" when "01100001", "10100110" when "01100010", "10100101" when "01100011", 
					"10101100" when "01100100", "10101111" when "01100101", "10101010" when "01100110", "10101001" when "01100111", 
					"10111000" when "01101000", "10111011" when "01101001", "10111110" when "01101010", "10111101" when "01101011", 
					"10110100" when "01101100", "10110111" when "01101101", "10110010" when "01101110", "10110001" when "01101111", 
					"10010000" when "01110000", "10010011" when "01110001", "10010110" when "01110010", "10010101" when "01110011", 
					"10011100" when "01110100", "10011111" when "01110101", "10011010" when "01110110", "10011001" when "01110111", 
					"10001000" when "01111000", "10001011" when "01111001", "10001110" when "01111010", "10001101" when "01111011", 
					"10000100" when "01111100", "10000111" when "01111101", "10000010" when "01111110", "10000001" when "01111111", 
					"11101001" when "10000000", "11101010" when "10000001", "11101111" when "10000010", "11101100" when "10000011", 
					"11100101" when "10000100", "11100110" when "10000101", "11100011" when "10000110", "11100000" when "10000111", 
					"11110001" when "10001000", "11110010" when "10001001", "11110111" when "10001010", "11110100" when "10001011", 
					"11111101" when "10001100", "11111110" when "10001101", "11111011" when "10001110", "11111000" when "10001111", 
					"11011001" when "10010000", "11011010" when "10010001", "11011111" when "10010010", "11011100" when "10010011", 
					"11010101" when "10010100", "11010110" when "10010101", "11010011" when "10010110", "11010000" when "10010111", 
					"11000001" when "10011000", "11000010" when "10011001", "11000111" when "10011010", "11000100" when "10011011", 
					"11001101" when "10011100", "11001110" when "10011101", "11001011" when "10011110", "11001000" when "10011111", 
					"10001001" when "10100000", "10001010" when "10100001", "10001111" when "10100010", "10001100" when "10100011", 
					"10000101" when "10100100", "10000110" when "10100101", "10000011" when "10100110", "10000000" when "10100111", 
					"10010001" when "10101000", "10010010" when "10101001", "10010111" when "10101010", "10010100" when "10101011", 
					"10011101" when "10101100", "10011110" when "10101101", "10011011" when "10101110", "10011000" when "10101111", 
					"10111001" when "10110000", "10111010" when "10110001", "10111111" when "10110010", "10111100" when "10110011", 
					"10110101" when "10110100", "10110110" when "10110101", "10110011" when "10110110", "10110000" when "10110111", 
					"10100001" when "10111000", "10100010" when "10111001", "10100111" when "10111010", "10100100" when "10111011", 
					"10101101" when "10111100", "10101110" when "10111101", "10101011" when "10111110", "10101000" when "10111111", 
					"00101001" when "11000000", "00101010" when "11000001", "00101111" when "11000010", "00101100" when "11000011", 
					"00100101" when "11000100", "00100110" when "11000101", "00100011" when "11000110", "00100000" when "11000111", 
					"00110001" when "11001000", "00110010" when "11001001", "00110111" when "11001010", "00110100" when "11001011", 
					"00111101" when "11001100", "00111110" when "11001101", "00111011" when "11001110", "00111000" when "11001111", 
					"00011001" when "11010000", "00011010" when "11010001", "00011111" when "11010010", "00011100" when "11010011", 
					"00010101" when "11010100", "00010110" when "11010101", "00010011" when "11010110", "00010000" when "11010111", 
					"00000001" when "11011000", "00000010" when "11011001", "00000111" when "11011010", "00000100" when "11011011", 
					"00001101" when "11011100", "00001110" when "11011101", "00001011" when "11011110", "00001000" when "11011111", 
					"01001001" when "11100000", "01001010" when "11100001", "01001111" when "11100010", "01001100" when "11100011", 
					"01000101" when "11100100", "01000110" when "11100101", "01000011" when "11100110", "01000000" when "11100111", 
					"01010001" when "11101000", "01010010" when "11101001", "01010111" when "11101010", "01010100" when "11101011", 
					"01011101" when "11101100", "01011110" when "11101101", "01011011" when "11101110", "01011000" when "11101111", 
					"01111001" when "11110000", "01111010" when "11110001", "01111111" when "11110010", "01111100" when "11110011", 
					"01110101" when "11110100", "01110110" when "11110101", "01110011" when "11110110", "01110000" when "11110111", 
					"01100001" when "11111000", "01100010" when "11111001", "01100111" when "11111010", "01100100" when "11111011", 
					"01101101" when "11111100", "01101110" when "11111101", "01101011" when "11111110", "01101000" when "11111111";

end mul_03_mem;

