----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:14:18 04/23/2021 
-- Design Name: 
-- Module Name:    mul_02_mem - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_02_mem is
	port (
			in_02 : in STD_LOGIC_VECTOR (7 downto 0);
			out_02 : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_02_mem;

architecture mul_02_mem of mul_02_mem is
begin

	with in_02 select
		out_02 <= "00000000" when "00000000", "00000010" when "00000001", "00000100" when "00000010", "00000110" when "00000011", 
					"00001000" when "00000100", "00001010" when "00000101", "00001100" when "00000110", "00001110" when "00000111", 
					"00010000" when "00001000", "00010010" when "00001001", "00010100" when "00001010", "00010110" when "00001011", 
					"00011000" when "00001100", "00011010" when "00001101", "00011100" when "00001110", "00011110" when "00001111", 
					"00100000" when "00010000", "00100010" when "00010001", "00100100" when "00010010", "00100110" when "00010011", 
					"00101000" when "00010100", "00101010" when "00010101", "00101100" when "00010110", "00101110" when "00010111", 
					"00110000" when "00011000", "00110010" when "00011001", "00110100" when "00011010", "00110110" when "00011011", 
					"00111000" when "00011100", "00111010" when "00011101", "00111100" when "00011110", "00111110" when "00011111", 
					"01000000" when "00100000", "01000010" when "00100001", "01000100" when "00100010", "01000110" when "00100011", 
					"01001000" when "00100100", "01001010" when "00100101", "01001100" when "00100110", "01001110" when "00100111", 
					"01010000" when "00101000", "01010010" when "00101001", "01010100" when "00101010", "01010110" when "00101011", 
					"01011000" when "00101100", "01011010" when "00101101", "01011100" when "00101110", "01011110" when "00101111", 
					"01100000" when "00110000", "01100010" when "00110001", "01100100" when "00110010", "01100110" when "00110011", 
					"01101000" when "00110100", "01101010" when "00110101", "01101100" when "00110110", "01101110" when "00110111", 
					"01110000" when "00111000", "01110010" when "00111001", "01110100" when "00111010", "01110110" when "00111011", 
					"01111000" when "00111100", "01111010" when "00111101", "01111100" when "00111110", "01111110" when "00111111", 
					"10000000" when "01000000", "10000010" when "01000001", "10000100" when "01000010", "10000110" when "01000011", 
					"10001000" when "01000100", "10001010" when "01000101", "10001100" when "01000110", "10001110" when "01000111", 
					"10010000" when "01001000", "10010010" when "01001001", "10010100" when "01001010", "10010110" when "01001011", 
					"10011000" when "01001100", "10011010" when "01001101", "10011100" when "01001110", "10011110" when "01001111", 
					"10100000" when "01010000", "10100010" when "01010001", "10100100" when "01010010", "10100110" when "01010011", 
					"10101000" when "01010100", "10101010" when "01010101", "10101100" when "01010110", "10101110" when "01010111", 
					"10110000" when "01011000", "10110010" when "01011001", "10110100" when "01011010", "10110110" when "01011011", 
					"10111000" when "01011100", "10111010" when "01011101", "10111100" when "01011110", "10111110" when "01011111", 
					"11000000" when "01100000", "11000010" when "01100001", "11000100" when "01100010", "11000110" when "01100011", 
					"11001000" when "01100100", "11001010" when "01100101", "11001100" when "01100110", "11001110" when "01100111", 
					"11010000" when "01101000", "11010010" when "01101001", "11010100" when "01101010", "11010110" when "01101011", 
					"11011000" when "01101100", "11011010" when "01101101", "11011100" when "01101110", "11011110" when "01101111", 
					"11100000" when "01110000", "11100010" when "01110001", "11100100" when "01110010", "11100110" when "01110011", 
					"11101000" when "01110100", "11101010" when "01110101", "11101100" when "01110110", "11101110" when "01110111", 
					"11110000" when "01111000", "11110010" when "01111001", "11110100" when "01111010", "11110110" when "01111011", 
					"11111000" when "01111100", "11111010" when "01111101", "11111100" when "01111110", "11111110" when "01111111", 
					"01101001" when "10000000", "01101011" when "10000001", "01101101" when "10000010", "01101111" when "10000011", 
					"01100001" when "10000100", "01100011" when "10000101", "01100101" when "10000110", "01100111" when "10000111", 
					"01111001" when "10001000", "01111011" when "10001001", "01111101" when "10001010", "01111111" when "10001011", 
					"01110001" when "10001100", "01110011" when "10001101", "01110101" when "10001110", "01110111" when "10001111", 
					"01001001" when "10010000", "01001011" when "10010001", "01001101" when "10010010", "01001111" when "10010011", 
					"01000001" when "10010100", "01000011" when "10010101", "01000101" when "10010110", "01000111" when "10010111", 
					"01011001" when "10011000", "01011011" when "10011001", "01011101" when "10011010", "01011111" when "10011011", 
					"01010001" when "10011100", "01010011" when "10011101", "01010101" when "10011110", "01010111" when "10011111", 
					"00101001" when "10100000", "00101011" when "10100001", "00101101" when "10100010", "00101111" when "10100011", 
					"00100001" when "10100100", "00100011" when "10100101", "00100101" when "10100110", "00100111" when "10100111", 
					"00111001" when "10101000", "00111011" when "10101001", "00111101" when "10101010", "00111111" when "10101011", 
					"00110001" when "10101100", "00110011" when "10101101", "00110101" when "10101110", "00110111" when "10101111", 
					"00001001" when "10110000", "00001011" when "10110001", "00001101" when "10110010", "00001111" when "10110011", 
					"00000001" when "10110100", "00000011" when "10110101", "00000101" when "10110110", "00000111" when "10110111", 
					"00011001" when "10111000", "00011011" when "10111001", "00011101" when "10111010", "00011111" when "10111011", 
					"00010001" when "10111100", "00010011" when "10111101", "00010101" when "10111110", "00010111" when "10111111", 
					"11101001" when "11000000", "11101011" when "11000001", "11101101" when "11000010", "11101111" when "11000011", 
					"11100001" when "11000100", "11100011" when "11000101", "11100101" when "11000110", "11100111" when "11000111", 
					"11111001" when "11001000", "11111011" when "11001001", "11111101" when "11001010", "11111111" when "11001011", 
					"11110001" when "11001100", "11110011" when "11001101", "11110101" when "11001110", "11110111" when "11001111", 
					"11001001" when "11010000", "11001011" when "11010001", "11001101" when "11010010", "11001111" when "11010011", 
					"11000001" when "11010100", "11000011" when "11010101", "11000101" when "11010110", "11000111" when "11010111", 
					"11011001" when "11011000", "11011011" when "11011001", "11011101" when "11011010", "11011111" when "11011011", 
					"11010001" when "11011100", "11010011" when "11011101", "11010101" when "11011110", "11010111" when "11011111", 
					"10101001" when "11100000", "10101011" when "11100001", "10101101" when "11100010", "10101111" when "11100011", 
					"10100001" when "11100100", "10100011" when "11100101", "10100101" when "11100110", "10100111" when "11100111", 
					"10111001" when "11101000", "10111011" when "11101001", "10111101" when "11101010", "10111111" when "11101011", 
					"10110001" when "11101100", "10110011" when "11101101", "10110101" when "11101110", "10110111" when "11101111", 
					"10001001" when "11110000", "10001011" when "11110001", "10001101" when "11110010", "10001111" when "11110011", 
					"10000001" when "11110100", "10000011" when "11110101", "10000101" when "11110110", "10000111" when "11110111", 
					"10011001" when "11111000", "10011011" when "11111001", "10011101" when "11111010", "10011111" when "11111011", 
					"10010001" when "11111100", "10010011" when "11111101", "10010101" when "11111110", "10010111" when "11111111";

end mul_02_mem;


