----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:47:46 04/21/2021 
-- Design Name: 
-- Module Name:    mult_5B_mem - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mult_5B_mem is
	port (
			in_5B : in STD_LOGIC_VECTOR (7 downto 0);
			out_5B : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mult_5B_mem;

architecture mult_5B_mem of mult_5B_mem is
begin

	with in_5B select
		out_5B <=	"00000000" when "00000000", "01011011" when "00000001", "10110110" when "00000010", "11101101" when "00000011",
					"00000101" when "00000100", "01011110" when "00000101", "10110011" when "00000110", "11101000" when "00000111",
					"00001010" when "00001000", "01010001" when "00001001", "10111100" when "00001010", "11100111" when "00001011",
					"00001111" when "00001100", "01010100" when "00001101", "10111001" when "00001110", "11100010" when "00001111",
					"00010100" when "00010000", "01001111" when "00010001", "10100010" when "00010010", "11111001" when "00010011",
					"00010001" when "00010100", "01001010" when "00010101", "10100111" when "00010110", "11111100" when "00010111",
					"00011110" when "00011000", "01000101" when "00011001", "10101000" when "00011010", "11110011" when "00011011",
					"00011011" when "00011100", "01000000" when "00011101", "10101101" when "00011110", "11110110" when "00011111",
					"00101000" when "00100000", "01110011" when "00100001", "10011110" when "00100010", "11000101" when "00100011",
					"00101101" when "00100100", "01110110" when "00100101", "10011011" when "00100110", "11000000" when "00100111",
					"00100010" when "00101000", "01111001" when "00101001", "10010100" when "00101010", "11001111" when "00101011",
					"00100111" when "00101100", "01111100" when "00101101", "10010001" when "00101110", "11001010" when "00101111",
					"00111100" when "00110000", "01100111" when "00110001", "10001010" when "00110010", "11010001" when "00110011",
					"00111001" when "00110100", "01100010" when "00110101", "10001111" when "00110110", "11010100" when "00110111",
					"00110110" when "00111000", "01101101" when "00111001", "10000000" when "00111010", "11011011" when "00111011",
					"00110011" when "00111100", "01101000" when "00111101", "10000101" when "00111110", "11011110" when "00111111",
					"01010000" when "01000000", "00001011" when "01000001", "11100110" when "01000010", "10111101" when "01000011",
					"01010101" when "01000100", "00001110" when "01000101", "11100011" when "01000110", "10111000" when "01000111",
					"01011010" when "01001000", "00000001" when "01001001", "11101100" when "01001010", "10110111" when "01001011",
					"01011111" when "01001100", "00000100" when "01001101", "11101001" when "01001110", "10110010" when "01001111",
					"01000100" when "01010000", "00011111" when "01010001", "11110010" when "01010010", "10101001" when "01010011",
					"01000001" when "01010100", "00011010" when "01010101", "11110111" when "01010110", "10101100" when "01010111",
					"01001110" when "01011000", "00010101" when "01011001", "11111000" when "01011010", "10100011" when "01011011",
					"01001011" when "01011100", "00010000" when "01011101", "11111101" when "01011110", "10100110" when "01011111",
					"01111000" when "01100000", "00100011" when "01100001", "11001110" when "01100010", "10010101" when "01100011",
					"01111101" when "01100100", "00100110" when "01100101", "11001011" when "01100110", "10010000" when "01100111",
					"01110010" when "01101000", "00101001" when "01101001", "11000100" when "01101010", "10011111" when "01101011",
					"01110111" when "01101100", "00101100" when "01101101", "11000001" when "01101110", "10011010" when "01101111",
					"01101100" when "01110000", "00110111" when "01110001", "11011010" when "01110010", "10000001" when "01110011",
					"01101001" when "01110100", "00110010" when "01110101", "11011111" when "01110110", "10000100" when "01110111",
					"01100110" when "01111000", "00111101" when "01111001", "11010000" when "01111010", "10001011" when "01111011",
					"01100011" when "01111100", "00111000" when "01111101", "11010101" when "01111110", "10001110" when "01111111",
					"10100000" when "10000000", "11111011" when "10000001", "00010110" when "10000010", "01001101" when "10000011",
					"10100101" when "10000100", "11111110" when "10000101", "00010011" when "10000110", "01001000" when "10000111",
					"10101010" when "10001000", "11110001" when "10001001", "00011100" when "10001010", "01000111" when "10001011",
					"10101111" when "10001100", "11110100" when "10001101", "00011001" when "10001110", "01000010" when "10001111",
					"10110100" when "10010000", "11101111" when "10010001", "00000010" when "10010010", "01011001" when "10010011",
					"10110001" when "10010100", "11101010" when "10010101", "00000111" when "10010110", "01011100" when "10010111",
					"10111110" when "10011000", "11100101" when "10011001", "00001000" when "10011010", "01010011" when "10011011",
					"10111011" when "10011100", "11100000" when "10011101", "00001101" when "10011110", "01010110" when "10011111",
					"10001000" when "10100000", "11010011" when "10100001", "00111110" when "10100010", "01100101" when "10100011",
					"10001101" when "10100100", "11010110" when "10100101", "00111011" when "10100110", "01100000" when "10100111",
					"10000010" when "10101000", "11011001" when "10101001", "00110100" when "10101010", "01101111" when "10101011",
					"10000111" when "10101100", "11011100" when "10101101", "00110001" when "10101110", "01101010" when "10101111",
					"10011100" when "10110000", "11000111" when "10110001", "00101010" when "10110010", "01110001" when "10110011",
					"10011001" when "10110100", "11000010" when "10110101", "00101111" when "10110110", "01110100" when "10110111",
					"10010110" when "10111000", "11001101" when "10111001", "00100000" when "10111010", "01111011" when "10111011",
					"10010011" when "10111100", "11001000" when "10111101", "00100101" when "10111110", "01111110" when "10111111",
					"11110000" when "11000000", "10101011" when "11000001", "01000110" when "11000010", "00011101" when "11000011",
					"11110101" when "11000100", "10101110" when "11000101", "01000011" when "11000110", "00011000" when "11000111",
					"11111010" when "11001000", "10100001" when "11001001", "01001100" when "11001010", "00010111" when "11001011",
					"11111111" when "11001100", "10100100" when "11001101", "01001001" when "11001110", "00010010" when "11001111",
					"11100100" when "11010000", "10111111" when "11010001", "01010010" when "11010010", "00001001" when "11010011",
					"11100001" when "11010100", "10111010" when "11010101", "01010111" when "11010110", "00001100" when "11010111",
					"11101110" when "11011000", "10110101" when "11011001", "01011000" when "11011010", "00000011" when "11011011",
					"11101011" when "11011100", "10110000" when "11011101", "01011101" when "11011110", "00000110" when "11011111",
					"11011000" when "11100000", "10000011" when "11100001", "01101110" when "11100010", "00110101" when "11100011",
					"11011101" when "11100100", "10000110" when "11100101", "01101011" when "11100110", "00110000" when "11100111",
					"11010010" when "11101000", "10001001" when "11101001", "01100100" when "11101010", "00111111" when "11101011",
					"11010111" when "11101100", "10001100" when "11101101", "01100001" when "11101110", "00111010" when "11101111",
					"11001100" when "11110000", "10010111" when "11110001", "01111010" when "11110010", "00100001" when "11110011",
					"11001001" when "11110100", "10010010" when "11110101", "01111111" when "11110110", "00100100" when "11110111",
					"11000110" when "11111000", "10011101" when "11111001", "01110000" when "11111010", "00101011" when "11111011",
					"11000011" when "11111100", "10011000" when "11111101", "01110101" when "11111110", "00101110" when "11111111";

end mult_5B_mem;