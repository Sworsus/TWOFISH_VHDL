----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:22:05 04/24/2021 
-- Design Name: 
-- Module Name:    mul_82_mem - mul_82_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_82_mem is
	port (
			in_82 : in STD_LOGIC_VECTOR (7 downto 0);
			out_82 : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_82_mem;

architecture mul_82_mem of mul_82_mem is

begin
	with in_82 select
	out_82 <= "00000000" when "00000000", 
				"10000010" when "00000001", 
				"01101101" when "00000010", 
				"11101111" when "00000011", 
				"11011010" when "00000100", 
				"01011000" when "00000101", 
				"10110111" when "00000110", 
				"00110101" when "00000111", 
				"11011101" when "00001000", 
				"01011111" when "00001001", 
				"10110000" when "00001010", 
				"00110010" when "00001011", 
				"00000111" when "00001100", 
				"10000101" when "00001101", 
				"01101010" when "00001110", 
				"11101000" when "00001111", 
				"11010011" when "00010000", 
				"01010001" when "00010001", 
				"10111110" when "00010010", 
				"00111100" when "00010011", 
				"00001001" when "00010100", 
				"10001011" when "00010101", 
				"01100100" when "00010110", 
				"11100110" when "00010111", 
				"00001110" when "00011000", 
				"10001100" when "00011001", 
				"01100011" when "00011010", 
				"11100001" when "00011011", 
				"11010100" when "00011100", 
				"01010110" when "00011101", 
				"10111001" when "00011110", 
				"00111011" when "00011111", 
				"11001111" when "00100000", 
				"01001101" when "00100001", 
				"10100010" when "00100010", 
				"00100000" when "00100011", 
				"00010101" when "00100100", 
				"10010111" when "00100101", 
				"01111000" when "00100110", 
				"11111010" when "00100111", 
				"00010010" when "00101000", 
				"10010000" when "00101001", 
				"01111111" when "00101010", 
				"11111101" when "00101011", 
				"11001000" when "00101100", 
				"01001010" when "00101101", 
				"10100101" when "00101110", 
				"00100111" when "00101111", 
				"00011100" when "00110000", 
				"10011110" when "00110001", 
				"01110001" when "00110010", 
				"11110011" when "00110011", 
				"11000110" when "00110100", 
				"01000100" when "00110101", 
				"10101011" when "00110110", 
				"00101001" when "00110111", 
				"11000001" when "00111000", 
				"01000011" when "00111001", 
				"10101100" when "00111010", 
				"00101110" when "00111011", 
				"00011011" when "00111100", 
				"10011001" when "00111101", 
				"01110110" when "00111110", 
				"11110100" when "00111111", 
				"11110111" when "01000000", 
				"01110101" when "01000001", 
				"10011010" when "01000010", 
				"00011000" when "01000011", 
				"00101101" when "01000100", 
				"10101111" when "01000101", 
				"01000000" when "01000110", 
				"11000010" when "01000111", 
				"00101010" when "01001000", 
				"10101000" when "01001001", 
				"01000111" when "01001010", 
				"11000101" when "01001011", 
				"11110000" when "01001100", 
				"01110010" when "01001101", 
				"10011101" when "01001110", 
				"00011111" when "01001111", 
				"00100100" when "01010000", 
				"10100110" when "01010001", 
				"01001001" when "01010010", 
				"11001011" when "01010011", 
				"11111110" when "01010100", 
				"01111100" when "01010101", 
				"10010011" when "01010110", 
				"00010001" when "01010111", 
				"11111001" when "01011000", 
				"01111011" when "01011001", 
				"10010100" when "01011010", 
				"00010110" when "01011011", 
				"00100011" when "01011100", 
				"10100001" when "01011101", 
				"01001110" when "01011110", 
				"11001100" when "01011111", 
				"00111000" when "01100000", 
				"10111010" when "01100001", 
				"01010101" when "01100010", 
				"11010111" when "01100011", 
				"11100010" when "01100100", 
				"01100000" when "01100101", 
				"10001111" when "01100110", 
				"00001101" when "01100111", 
				"11100101" when "01101000", 
				"01100111" when "01101001", 
				"10001000" when "01101010", 
				"00001010" when "01101011", 
				"00111111" when "01101100", 
				"10111101" when "01101101", 
				"01010010" when "01101110", 
				"11010000" when "01101111", 
				"11101011" when "01110000", 
				"01101001" when "01110001", 
				"10000110" when "01110010", 
				"00000100" when "01110011", 
				"00110001" when "01110100", 
				"10110011" when "01110101", 
				"01011100" when "01110110", 
				"11011110" when "01110111", 
				"00110110" when "01111000", 
				"10110100" when "01111001", 
				"01011011" when "01111010", 
				"11011001" when "01111011", 
				"11101100" when "01111100", 
				"01101110" when "01111101", 
				"10000001" when "01111110", 
				"00000011" when "01111111", 
				"10000111" when "10000000", 
				"00000101" when "10000001", 
				"11101010" when "10000010", 
				"01101000" when "10000011", 
				"01011101" when "10000100", 
				"11011111" when "10000101", 
				"00110000" when "10000110", 
				"10110010" when "10000111", 
				"01011010" when "10001000", 
				"11011000" when "10001001", 
				"00110111" when "10001010", 
				"10110101" when "10001011", 
				"10000000" when "10001100", 
				"00000010" when "10001101", 
				"11101101" when "10001110", 
				"01101111" when "10001111", 
				"01010100" when "10010000", 
				"11010110" when "10010001", 
				"00111001" when "10010010", 
				"10111011" when "10010011", 
				"10001110" when "10010100", 
				"00001100" when "10010101", 
				"11100011" when "10010110", 
				"01100001" when "10010111", 
				"10001001" when "10011000", 
				"00001011" when "10011001", 
				"11100100" when "10011010", 
				"01100110" when "10011011", 
				"01010011" when "10011100", 
				"11010001" when "10011101", 
				"00111110" when "10011110", 
				"10111100" when "10011111", 
				"01001000" when "10100000", 
				"11001010" when "10100001", 
				"00100101" when "10100010", 
				"10100111" when "10100011", 
				"10010010" when "10100100", 
				"00010000" when "10100101", 
				"11111111" when "10100110", 
				"01111101" when "10100111", 
				"10010101" when "10101000", 
				"00010111" when "10101001", 
				"11111000" when "10101010", 
				"01111010" when "10101011", 
				"01001111" when "10101100", 
				"11001101" when "10101101", 
				"00100010" when "10101110", 
				"10100000" when "10101111", 
				"10011011" when "10110000", 
				"00011001" when "10110001", 
				"11110110" when "10110010", 
				"01110100" when "10110011", 
				"01000001" when "10110100", 
				"11000011" when "10110101", 
				"00101100" when "10110110", 
				"10101110" when "10110111", 
				"01000110" when "10111000", 
				"11000100" when "10111001", 
				"00101011" when "10111010", 
				"10101001" when "10111011", 
				"10011100" when "10111100", 
				"00011110" when "10111101", 
				"11110001" when "10111110", 
				"01110011" when "10111111", 
				"01110000" when "11000000", 
				"11110010" when "11000001", 
				"00011101" when "11000010", 
				"10011111" when "11000011", 
				"10101010" when "11000100", 
				"00101000" when "11000101", 
				"11000111" when "11000110", 
				"01000101" when "11000111", 
				"10101101" when "11001000", 
				"00101111" when "11001001", 
				"11000000" when "11001010", 
				"01000010" when "11001011", 
				"01110111" when "11001100", 
				"11110101" when "11001101", 
				"00011010" when "11001110", 
				"10011000" when "11001111", 
				"10100011" when "11010000", 
				"00100001" when "11010001", 
				"11001110" when "11010010", 
				"01001100" when "11010011", 
				"01111001" when "11010100", 
				"11111011" when "11010101", 
				"00010100" when "11010110", 
				"10010110" when "11010111", 
				"01111110" when "11011000", 
				"11111100" when "11011001", 
				"00010011" when "11011010", 
				"10010001" when "11011011", 
				"10100100" when "11011100", 
				"00100110" when "11011101", 
				"11001001" when "11011110", 
				"01001011" when "11011111", 
				"10111111" when "11100000", 
				"00111101" when "11100001", 
				"11010010" when "11100010", 
				"01010000" when "11100011", 
				"01100101" when "11100100", 
				"11100111" when "11100101", 
				"00001000" when "11100110", 
				"10001010" when "11100111", 
				"01100010" when "11101000", 
				"11100000" when "11101001", 
				"00001111" when "11101010", 
				"10001101" when "11101011", 
				"10111000" when "11101100", 
				"00111010" when "11101101", 
				"11010101" when "11101110", 
				"01010111" when "11101111", 
				"01101100" when "11110000", 
				"11101110" when "11110001", 
				"00000001" when "11110010", 
				"10000011" when "11110011", 
				"10110110" when "11110100", 
				"00110100" when "11110101", 
				"11011011" when "11110110", 
				"01011001" when "11110111", 
				"10110001" when "11111000", 
				"00110011" when "11111001", 
				"11011100" when "11111010", 
				"01011110" when "11111011", 
				"01101011" when "11111100", 
				"11101001" when "11111101", 
				"00000110" when "11111110", 
				"10000100" when "11111111";

end mul_82_mem;

