----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    01:08:32 04/24/2021 
-- Design Name: 
-- Module Name:    mul_56_mem - mul_56_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_56_mem is
	port (
			in_56 : in STD_LOGIC_VECTOR (7 downto 0);
			out_56 : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_56_mem;

architecture mul_56_mem of mul_56_mem is
begin
	
	with in_56 select
	out_56 <= "00000000" when "00000000", 
				"01010110" when "00000001", 
				"10101100" when "00000010", 
				"11111010" when "00000011", 
				"00110001" when "00000100", 
				"01100111" when "00000101", 
				"10011101" when "00000110", 
				"11001011" when "00000111", 
				"01100010" when "00001000", 
				"00110100" when "00001001", 
				"11001110" when "00001010", 
				"10011000" when "00001011", 
				"01010011" when "00001100", 
				"00000101" when "00001101", 
				"11111111" when "00001110", 
				"10101001" when "00001111", 
				"11000100" when "00010000", 
				"10010010" when "00010001", 
				"01101000" when "00010010", 
				"00111110" when "00010011", 
				"11110101" when "00010100", 
				"10100011" when "00010101", 
				"01011001" when "00010110", 
				"00001111" when "00010111", 
				"10100110" when "00011000", 
				"11110000" when "00011001", 
				"00001010" when "00011010", 
				"01011100" when "00011011", 
				"10010111" when "00011100", 
				"11000001" when "00011101", 
				"00111011" when "00011110", 
				"01101101" when "00011111", 
				"11100001" when "00100000", 
				"10110111" when "00100001", 
				"01001101" when "00100010", 
				"00011011" when "00100011", 
				"11010000" when "00100100", 
				"10000110" when "00100101", 
				"01111100" when "00100110", 
				"00101010" when "00100111", 
				"10000011" when "00101000", 
				"11010101" when "00101001", 
				"00101111" when "00101010", 
				"01111001" when "00101011", 
				"10110010" when "00101100", 
				"11100100" when "00101101", 
				"00011110" when "00101110", 
				"01001000" when "00101111", 
				"00100101" when "00110000", 
				"01110011" when "00110001", 
				"10001001" when "00110010", 
				"11011111" when "00110011", 
				"00010100" when "00110100", 
				"01000010" when "00110101", 
				"10111000" when "00110110", 
				"11101110" when "00110111", 
				"01000111" when "00111000", 
				"00010001" when "00111001", 
				"11101011" when "00111010", 
				"10111101" when "00111011", 
				"01110110" when "00111100", 
				"00100000" when "00111101", 
				"11011010" when "00111110", 
				"10001100" when "00111111", 
				"10101011" when "01000000", 
				"11111101" when "01000001", 
				"00000111" when "01000010", 
				"01010001" when "01000011", 
				"10011010" when "01000100", 
				"11001100" when "01000101", 
				"00110110" when "01000110", 
				"01100000" when "01000111", 
				"11001001" when "01001000", 
				"10011111" when "01001001", 
				"01100101" when "01001010", 
				"00110011" when "01001011", 
				"11111000" when "01001100", 
				"10101110" when "01001101", 
				"01010100" when "01001110", 
				"00000010" when "01001111", 
				"01101111" when "01010000", 
				"00111001" when "01010001", 
				"11000011" when "01010010", 
				"10010101" when "01010011", 
				"01011110" when "01010100", 
				"00001000" when "01010101", 
				"11110010" when "01010110", 
				"10100100" when "01010111", 
				"00001101" when "01011000", 
				"01011011" when "01011001", 
				"10100001" when "01011010", 
				"11110111" when "01011011", 
				"00111100" when "01011100", 
				"01101010" when "01011101", 
				"10010000" when "01011110", 
				"11000110" when "01011111", 
				"01001010" when "01100000", 
				"00011100" when "01100001", 
				"11100110" when "01100010", 
				"10110000" when "01100011", 
				"01111011" when "01100100", 
				"00101101" when "01100101", 
				"11010111" when "01100110", 
				"10000001" when "01100111", 
				"00101000" when "01101000", 
				"01111110" when "01101001", 
				"10000100" when "01101010", 
				"11010010" when "01101011", 
				"00011001" when "01101100", 
				"01001111" when "01101101", 
				"10110101" when "01101110", 
				"11100011" when "01101111", 
				"10001110" when "01110000", 
				"11011000" when "01110001", 
				"00100010" when "01110010", 
				"01110100" when "01110011", 
				"10111111" when "01110100", 
				"11101001" when "01110101", 
				"00010011" when "01110110", 
				"01000101" when "01110111", 
				"11101100" when "01111000", 
				"10111010" when "01111001", 
				"01000000" when "01111010", 
				"00010110" when "01111011", 
				"11011101" when "01111100", 
				"10001011" when "01111101", 
				"01110001" when "01111110", 
				"00100111" when "01111111", 
				"00111111" when "10000000", 
				"01101001" when "10000001", 
				"10010011" when "10000010", 
				"11000101" when "10000011", 
				"00001110" when "10000100", 
				"01011000" when "10000101", 
				"10100010" when "10000110", 
				"11110100" when "10000111", 
				"01011101" when "10001000", 
				"00001011" when "10001001", 
				"11110001" when "10001010", 
				"10100111" when "10001011", 
				"01101100" when "10001100", 
				"00111010" when "10001101", 
				"11000000" when "10001110", 
				"10010110" when "10001111", 
				"11111011" when "10010000", 
				"10101101" when "10010001", 
				"01010111" when "10010010", 
				"00000001" when "10010011", 
				"11001010" when "10010100", 
				"10011100" when "10010101", 
				"01100110" when "10010110", 
				"00110000" when "10010111", 
				"10011001" when "10011000", 
				"11001111" when "10011001", 
				"00110101" when "10011010", 
				"01100011" when "10011011", 
				"10101000" when "10011100", 
				"11111110" when "10011101", 
				"00000100" when "10011110", 
				"01010010" when "10011111", 
				"11011110" when "10100000", 
				"10001000" when "10100001", 
				"01110010" when "10100010", 
				"00100100" when "10100011", 
				"11101111" when "10100100", 
				"10111001" when "10100101", 
				"01000011" when "10100110", 
				"00010101" when "10100111", 
				"10111100" when "10101000", 
				"11101010" when "10101001", 
				"00010000" when "10101010", 
				"01000110" when "10101011", 
				"10001101" when "10101100", 
				"11011011" when "10101101", 
				"00100001" when "10101110", 
				"01110111" when "10101111", 
				"00011010" when "10110000", 
				"01001100" when "10110001", 
				"10110110" when "10110010", 
				"11100000" when "10110011", 
				"00101011" when "10110100", 
				"01111101" when "10110101", 
				"10000111" when "10110110", 
				"11010001" when "10110111", 
				"01111000" when "10111000", 
				"00101110" when "10111001", 
				"11010100" when "10111010", 
				"10000010" when "10111011", 
				"01001001" when "10111100", 
				"00011111" when "10111101", 
				"11100101" when "10111110", 
				"10110011" when "10111111", 
				"10010100" when "11000000", 
				"11000010" when "11000001", 
				"00111000" when "11000010", 
				"01101110" when "11000011", 
				"10100101" when "11000100", 
				"11110011" when "11000101", 
				"00001001" when "11000110", 
				"01011111" when "11000111", 
				"11110110" when "11001000", 
				"10100000" when "11001001", 
				"01011010" when "11001010", 
				"00001100" when "11001011", 
				"11000111" when "11001100", 
				"10010001" when "11001101", 
				"01101011" when "11001110", 
				"00111101" when "11001111", 
				"01010000" when "11010000", 
				"00000110" when "11010001", 
				"11111100" when "11010010", 
				"10101010" when "11010011", 
				"01100001" when "11010100", 
				"00110111" when "11010101", 
				"11001101" when "11010110", 
				"10011011" when "11010111", 
				"00110010" when "11011000", 
				"01100100" when "11011001", 
				"10011110" when "11011010", 
				"11001000" when "11011011", 
				"00000011" when "11011100", 
				"01010101" when "11011101", 
				"10101111" when "11011110", 
				"11111001" when "11011111", 
				"01110101" when "11100000", 
				"00100011" when "11100001", 
				"11011001" when "11100010", 
				"10001111" when "11100011", 
				"01000100" when "11100100", 
				"00010010" when "11100101", 
				"11101000" when "11100110", 
				"10111110" when "11100111", 
				"00010111" when "11101000", 
				"01000001" when "11101001", 
				"10111011" when "11101010", 
				"11101101" when "11101011", 
				"00100110" when "11101100", 
				"01110000" when "11101101", 
				"10001010" when "11101110", 
				"11011100" when "11101111", 
				"10110001" when "11110000", 
				"11100111" when "11110001", 
				"00011101" when "11110010", 
				"01001011" when "11110011", 
				"10000000" when "11110100", 
				"11010110" when "11110101", 
				"00101100" when "11110110", 
				"01111010" when "11110111", 
				"11010011" when "11111000", 
				"10000101" when "11111001", 
				"01111111" when "11111010", 
				"00101001" when "11111011", 
				"11100010" when "11111100", 
				"10110100" when "11111101", 
				"01001110" when "11111110", 
				"00011000" when "11111111";

end mul_56_mem;

