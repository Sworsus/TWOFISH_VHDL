----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    01:41:22 04/24/2021 
-- Design Name: 
-- Module Name:    mul_5A_mem - mul_5A_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_5A_mem is
	port (
			in_5A : in STD_LOGIC_VECTOR (7 downto 0);
			out_5A : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_5A_mem;

architecture mul_5A_mem of mul_5A_mem is

begin

	with in_5A select
	out_5A <= "00000000" when "00000000", 
				"01011010" when "00000001", 
				"10110100" when "00000010", 
				"11101110" when "00000011", 
				"00000001" when "00000100", 
				"01011011" when "00000101", 
				"10110101" when "00000110", 
				"11101111" when "00000111", 
				"00000010" when "00001000", 
				"01011000" when "00001001", 
				"10110110" when "00001010", 
				"11101100" when "00001011", 
				"00000011" when "00001100", 
				"01011001" when "00001101", 
				"10110111" when "00001110", 
				"11101101" when "00001111", 
				"00000100" when "00010000", 
				"01011110" when "00010001", 
				"10110000" when "00010010", 
				"11101010" when "00010011", 
				"00000101" when "00010100", 
				"01011111" when "00010101", 
				"10110001" when "00010110", 
				"11101011" when "00010111", 
				"00000110" when "00011000", 
				"01011100" when "00011001", 
				"10110010" when "00011010", 
				"11101000" when "00011011", 
				"00000111" when "00011100", 
				"01011101" when "00011101", 
				"10110011" when "00011110", 
				"11101001" when "00011111", 
				"00001000" when "00100000", 
				"01010010" when "00100001", 
				"10111100" when "00100010", 
				"11100110" when "00100011", 
				"00001001" when "00100100", 
				"01010011" when "00100101", 
				"10111101" when "00100110", 
				"11100111" when "00100111", 
				"00001010" when "00101000", 
				"01010000" when "00101001", 
				"10111110" when "00101010", 
				"11100100" when "00101011", 
				"00001011" when "00101100", 
				"01010001" when "00101101", 
				"10111111" when "00101110", 
				"11100101" when "00101111", 
				"00001100" when "00110000", 
				"01010110" when "00110001", 
				"10111000" when "00110010", 
				"11100010" when "00110011", 
				"00001101" when "00110100", 
				"01010111" when "00110101", 
				"10111001" when "00110110", 
				"11100011" when "00110111", 
				"00001110" when "00111000", 
				"01010100" when "00111001", 
				"10111010" when "00111010", 
				"11100000" when "00111011", 
				"00001111" when "00111100", 
				"01010101" when "00111101", 
				"10111011" when "00111110", 
				"11100001" when "00111111", 
				"00010000" when "01000000", 
				"01001010" when "01000001", 
				"10100100" when "01000010", 
				"11111110" when "01000011", 
				"00010001" when "01000100", 
				"01001011" when "01000101", 
				"10100101" when "01000110", 
				"11111111" when "01000111", 
				"00010010" when "01001000", 
				"01001000" when "01001001", 
				"10100110" when "01001010", 
				"11111100" when "01001011", 
				"00010011" when "01001100", 
				"01001001" when "01001101", 
				"10100111" when "01001110", 
				"11111101" when "01001111", 
				"00010100" when "01010000", 
				"01001110" when "01010001", 
				"10100000" when "01010010", 
				"11111010" when "01010011", 
				"00010101" when "01010100", 
				"01001111" when "01010101", 
				"10100001" when "01010110", 
				"11111011" when "01010111", 
				"00010110" when "01011000", 
				"01001100" when "01011001", 
				"10100010" when "01011010", 
				"11111000" when "01011011", 
				"00010111" when "01011100", 
				"01001101" when "01011101", 
				"10100011" when "01011110", 
				"11111001" when "01011111", 
				"00011000" when "01100000", 
				"01000010" when "01100001", 
				"10101100" when "01100010", 
				"11110110" when "01100011", 
				"00011001" when "01100100", 
				"01000011" when "01100101", 
				"10101101" when "01100110", 
				"11110111" when "01100111", 
				"00011010" when "01101000", 
				"01000000" when "01101001", 
				"10101110" when "01101010", 
				"11110100" when "01101011", 
				"00011011" when "01101100", 
				"01000001" when "01101101", 
				"10101111" when "01101110", 
				"11110101" when "01101111", 
				"00011100" when "01110000", 
				"01000110" when "01110001", 
				"10101000" when "01110010", 
				"11110010" when "01110011", 
				"00011101" when "01110100", 
				"01000111" when "01110101", 
				"10101001" when "01110110", 
				"11110011" when "01110111", 
				"00011110" when "01111000", 
				"01000100" when "01111001", 
				"10101010" when "01111010", 
				"11110000" when "01111011", 
				"00011111" when "01111100", 
				"01000101" when "01111101", 
				"10101011" when "01111110", 
				"11110001" when "01111111", 
				"00100000" when "10000000", 
				"01111010" when "10000001", 
				"10010100" when "10000010", 
				"11001110" when "10000011", 
				"00100001" when "10000100", 
				"01111011" when "10000101", 
				"10010101" when "10000110", 
				"11001111" when "10000111", 
				"00100010" when "10001000", 
				"01111000" when "10001001", 
				"10010110" when "10001010", 
				"11001100" when "10001011", 
				"00100011" when "10001100", 
				"01111001" when "10001101", 
				"10010111" when "10001110", 
				"11001101" when "10001111", 
				"00100100" when "10010000", 
				"01111110" when "10010001", 
				"10010000" when "10010010", 
				"11001010" when "10010011", 
				"00100101" when "10010100", 
				"01111111" when "10010101", 
				"10010001" when "10010110", 
				"11001011" when "10010111", 
				"00100110" when "10011000", 
				"01111100" when "10011001", 
				"10010010" when "10011010", 
				"11001000" when "10011011", 
				"00100111" when "10011100", 
				"01111101" when "10011101", 
				"10010011" when "10011110", 
				"11001001" when "10011111", 
				"00101000" when "10100000", 
				"01110010" when "10100001", 
				"10011100" when "10100010", 
				"11000110" when "10100011", 
				"00101001" when "10100100", 
				"01110011" when "10100101", 
				"10011101" when "10100110", 
				"11000111" when "10100111", 
				"00101010" when "10101000", 
				"01110000" when "10101001", 
				"10011110" when "10101010", 
				"11000100" when "10101011", 
				"00101011" when "10101100", 
				"01110001" when "10101101", 
				"10011111" when "10101110", 
				"11000101" when "10101111", 
				"00101100" when "10110000", 
				"01110110" when "10110001", 
				"10011000" when "10110010", 
				"11000010" when "10110011", 
				"00101101" when "10110100", 
				"01110111" when "10110101", 
				"10011001" when "10110110", 
				"11000011" when "10110111", 
				"00101110" when "10111000", 
				"01110100" when "10111001", 
				"10011010" when "10111010", 
				"11000000" when "10111011", 
				"00101111" when "10111100", 
				"01110101" when "10111101", 
				"10011011" when "10111110", 
				"11000001" when "10111111", 
				"00110000" when "11000000", 
				"01101010" when "11000001", 
				"10000100" when "11000010", 
				"11011110" when "11000011", 
				"00110001" when "11000100", 
				"01101011" when "11000101", 
				"10000101" when "11000110", 
				"11011111" when "11000111", 
				"00110010" when "11001000", 
				"01101000" when "11001001", 
				"10000110" when "11001010", 
				"11011100" when "11001011", 
				"00110011" when "11001100", 
				"01101001" when "11001101", 
				"10000111" when "11001110", 
				"11011101" when "11001111", 
				"00110100" when "11010000", 
				"01101110" when "11010001", 
				"10000000" when "11010010", 
				"11011010" when "11010011", 
				"00110101" when "11010100", 
				"01101111" when "11010101", 
				"10000001" when "11010110", 
				"11011011" when "11010111", 
				"00110110" when "11011000", 
				"01101100" when "11011001", 
				"10000010" when "11011010", 
				"11011000" when "11011011", 
				"00110111" when "11011100", 
				"01101101" when "11011101", 
				"10000011" when "11011110", 
				"11011001" when "11011111", 
				"00111000" when "11100000", 
				"01100010" when "11100001", 
				"10001100" when "11100010", 
				"11010110" when "11100011", 
				"00111001" when "11100100", 
				"01100011" when "11100101", 
				"10001101" when "11100110", 
				"11010111" when "11100111", 
				"00111010" when "11101000", 
				"01100000" when "11101001", 
				"10001110" when "11101010", 
				"11010100" when "11101011", 
				"00111011" when "11101100", 
				"01100001" when "11101101", 
				"10001111" when "11101110", 
				"11010101" when "11101111", 
				"00111100" when "11110000", 
				"01100110" when "11110001", 
				"10001000" when "11110010", 
				"11010010" when "11110011", 
				"00111101" when "11110100", 
				"01100111" when "11110101", 
				"10001001" when "11110110", 
				"11010011" when "11110111", 
				"00111110" when "11111000", 
				"01100100" when "11111001", 
				"10001010" when "11111010", 
				"11010000" when "11111011", 
				"00111111" when "11111100", 
				"01100101" when "11111101", 
				"10001011" when "11111110", 
				"11010001" when "11111111";

end mul_5A_mem;

