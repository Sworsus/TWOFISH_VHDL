----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:54:49 04/24/2021 
-- Design Name: 
-- Module Name:    mul_DB_mem - mul_DB_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_DB_mem is
	port (
			in_DB : in STD_LOGIC_VECTOR (7 downto 0);
			out_DB : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_DB_mem;

architecture mul_DB_mem of mul_DB_mem is

begin

	with in_DB select
	out_DB <= "00000000" when "00000000", 
				"11011011" when "00000001", 
				"11011111" when "00000010", 
				"00000100" when "00000011", 
				"11010111" when "00000100", 
				"00001100" when "00000101", 
				"00001000" when "00000110", 
				"11010011" when "00000111", 
				"11000111" when "00001000", 
				"00011100" when "00001001", 
				"00011000" when "00001010", 
				"11000011" when "00001011", 
				"00010000" when "00001100", 
				"11001011" when "00001101", 
				"11001111" when "00001110", 
				"00010100" when "00001111", 
				"11100111" when "00010000", 
				"00111100" when "00010001", 
				"00111000" when "00010010", 
				"11100011" when "00010011", 
				"00110000" when "00010100", 
				"11101011" when "00010101", 
				"11101111" when "00010110", 
				"00110100" when "00010111", 
				"00100000" when "00011000", 
				"11111011" when "00011001", 
				"11111111" when "00011010", 
				"00100100" when "00011011", 
				"11110111" when "00011100", 
				"00101100" when "00011101", 
				"00101000" when "00011110", 
				"11110011" when "00011111", 
				"10100111" when "00100000", 
				"01111100" when "00100001", 
				"01111000" when "00100010", 
				"10100011" when "00100011", 
				"01110000" when "00100100", 
				"10101011" when "00100101", 
				"10101111" when "00100110", 
				"01110100" when "00100111", 
				"01100000" when "00101000", 
				"10111011" when "00101001", 
				"10111111" when "00101010", 
				"01100100" when "00101011", 
				"10110111" when "00101100", 
				"01101100" when "00101101", 
				"01101000" when "00101110", 
				"10110011" when "00101111", 
				"01000000" when "00110000", 
				"10011011" when "00110001", 
				"10011111" when "00110010", 
				"01000100" when "00110011", 
				"10010111" when "00110100", 
				"01001100" when "00110101", 
				"01001000" when "00110110", 
				"10010011" when "00110111", 
				"10000111" when "00111000", 
				"01011100" when "00111001", 
				"01011000" when "00111010", 
				"10000011" when "00111011", 
				"01010000" when "00111100", 
				"10001011" when "00111101", 
				"10001111" when "00111110", 
				"01010100" when "00111111", 
				"00100111" when "01000000", 
				"11111100" when "01000001", 
				"11111000" when "01000010", 
				"00100011" when "01000011", 
				"11110000" when "01000100", 
				"00101011" when "01000101", 
				"00101111" when "01000110", 
				"11110100" when "01000111", 
				"11100000" when "01001000", 
				"00111011" when "01001001", 
				"00111111" when "01001010", 
				"11100100" when "01001011", 
				"00110111" when "01001100", 
				"11101100" when "01001101", 
				"11101000" when "01001110", 
				"00110011" when "01001111", 
				"11000000" when "01010000", 
				"00011011" when "01010001", 
				"00011111" when "01010010", 
				"11000100" when "01010011", 
				"00010111" when "01010100", 
				"11001100" when "01010101", 
				"11001000" when "01010110", 
				"00010011" when "01010111", 
				"00000111" when "01011000", 
				"11011100" when "01011001", 
				"11011000" when "01011010", 
				"00000011" when "01011011", 
				"11010000" when "01011100", 
				"00001011" when "01011101", 
				"00001111" when "01011110", 
				"11010100" when "01011111", 
				"10000000" when "01100000", 
				"01011011" when "01100001", 
				"01011111" when "01100010", 
				"10000100" when "01100011", 
				"01010111" when "01100100", 
				"10001100" when "01100101", 
				"10001000" when "01100110", 
				"01010011" when "01100111", 
				"01000111" when "01101000", 
				"10011100" when "01101001", 
				"10011000" when "01101010", 
				"01000011" when "01101011", 
				"10010000" when "01101100", 
				"01001011" when "01101101", 
				"01001111" when "01101110", 
				"10010100" when "01101111", 
				"01100111" when "01110000", 
				"10111100" when "01110001", 
				"10111000" when "01110010", 
				"01100011" when "01110011", 
				"10110000" when "01110100", 
				"01101011" when "01110101", 
				"01101111" when "01110110", 
				"10110100" when "01110111", 
				"10100000" when "01111000", 
				"01111011" when "01111001", 
				"01111111" when "01111010", 
				"10100100" when "01111011", 
				"01110111" when "01111100", 
				"10101100" when "01111101", 
				"10101000" when "01111110", 
				"01110011" when "01111111", 
				"01001110" when "10000000", 
				"10010101" when "10000001", 
				"10010001" when "10000010", 
				"01001010" when "10000011", 
				"10011001" when "10000100", 
				"01000010" when "10000101", 
				"01000110" when "10000110", 
				"10011101" when "10000111", 
				"10001001" when "10001000", 
				"01010010" when "10001001", 
				"01010110" when "10001010", 
				"10001101" when "10001011", 
				"01011110" when "10001100", 
				"10000101" when "10001101", 
				"10000001" when "10001110", 
				"01011010" when "10001111", 
				"10101001" when "10010000", 
				"01110010" when "10010001", 
				"01110110" when "10010010", 
				"10101101" when "10010011", 
				"01111110" when "10010100", 
				"10100101" when "10010101", 
				"10100001" when "10010110", 
				"01111010" when "10010111", 
				"01101110" when "10011000", 
				"10110101" when "10011001", 
				"10110001" when "10011010", 
				"01101010" when "10011011", 
				"10111001" when "10011100", 
				"01100010" when "10011101", 
				"01100110" when "10011110", 
				"10111101" when "10011111", 
				"11101001" when "10100000", 
				"00110010" when "10100001", 
				"00110110" when "10100010", 
				"11101101" when "10100011", 
				"00111110" when "10100100", 
				"11100101" when "10100101", 
				"11100001" when "10100110", 
				"00111010" when "10100111", 
				"00101110" when "10101000", 
				"11110101" when "10101001", 
				"11110001" when "10101010", 
				"00101010" when "10101011", 
				"11111001" when "10101100", 
				"00100010" when "10101101", 
				"00100110" when "10101110", 
				"11111101" when "10101111", 
				"00001110" when "10110000", 
				"11010101" when "10110001", 
				"11010001" when "10110010", 
				"00001010" when "10110011", 
				"11011001" when "10110100", 
				"00000010" when "10110101", 
				"00000110" when "10110110", 
				"11011101" when "10110111", 
				"11001001" when "10111000", 
				"00010010" when "10111001", 
				"00010110" when "10111010", 
				"11001101" when "10111011", 
				"00011110" when "10111100", 
				"11000101" when "10111101", 
				"11000001" when "10111110", 
				"00011010" when "10111111", 
				"01101001" when "11000000", 
				"10110010" when "11000001", 
				"10110110" when "11000010", 
				"01101101" when "11000011", 
				"10111110" when "11000100", 
				"01100101" when "11000101", 
				"01100001" when "11000110", 
				"10111010" when "11000111", 
				"10101110" when "11001000", 
				"01110101" when "11001001", 
				"01110001" when "11001010", 
				"10101010" when "11001011", 
				"01111001" when "11001100", 
				"10100010" when "11001101", 
				"10100110" when "11001110", 
				"01111101" when "11001111", 
				"10001110" when "11010000", 
				"01010101" when "11010001", 
				"01010001" when "11010010", 
				"10001010" when "11010011", 
				"01011001" when "11010100", 
				"10000010" when "11010101", 
				"10000110" when "11010110", 
				"01011101" when "11010111", 
				"01001001" when "11011000", 
				"10010010" when "11011001", 
				"10010110" when "11011010", 
				"01001101" when "11011011", 
				"10011110" when "11011100", 
				"01000101" when "11011101", 
				"01000001" when "11011110", 
				"10011010" when "11011111", 
				"11001110" when "11100000", 
				"00010101" when "11100001", 
				"00010001" when "11100010", 
				"11001010" when "11100011", 
				"00011001" when "11100100", 
				"11000010" when "11100101", 
				"11000110" when "11100110", 
				"00011101" when "11100111", 
				"00001001" when "11101000", 
				"11010010" when "11101001", 
				"11010110" when "11101010", 
				"00001101" when "11101011", 
				"11011110" when "11101100", 
				"00000101" when "11101101", 
				"00000001" when "11101110", 
				"11011010" when "11101111", 
				"00101001" when "11110000", 
				"11110010" when "11110001", 
				"11110110" when "11110010", 
				"00101101" when "11110011", 
				"11111110" when "11110100", 
				"00100101" when "11110101", 
				"00100001" when "11110110", 
				"11111010" when "11110111", 
				"11101110" when "11111000", 
				"00110101" when "11111001", 
				"00110001" when "11111010", 
				"11101010" when "11111011", 
				"00111001" when "11111100", 
				"11100010" when "11111101", 
				"11100110" when "11111110", 
				"00111101" when "11111111";

end mul_DB_mem;

