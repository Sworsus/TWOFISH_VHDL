----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:04:44 04/23/2021 
-- Design Name: 
-- Module Name:    mul_1E_mem - mul_1E_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_1E_mem is
	port (
			in_1E : in STD_LOGIC_VECTOR (7 downto 0);
			out_1E : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_1E_mem;

architecture mul_1E_mem of mul_1E_mem is

begin

		with in_1E select
			out_1E <= "00000000" when "00000000", 
						"00011110" when "00000001", 
						"00111100" when "00000010", 
						"00100010" when "00000011", 
						"01111000" when "00000100", 
						"01100110" when "00000101", 
						"01000100" when "00000110", 
						"01011010" when "00000111", 
						"11110000" when "00001000", 
						"11101110" when "00001001", 
						"11001100" when "00001010", 
						"11010010" when "00001011", 
						"10001000" when "00001100", 
						"10010110" when "00001101", 
						"10110100" when "00001110", 
						"10101010" when "00001111", 
						"10001001" when "00010000", 
						"10010111" when "00010001", 
						"10110101" when "00010010", 
						"10101011" when "00010011", 
						"11110001" when "00010100", 
						"11101111" when "00010101", 
						"11001101" when "00010110", 
						"11010011" when "00010111", 
						"01111001" when "00011000", 
						"01100111" when "00011001", 
						"01000101" when "00011010", 
						"01011011" when "00011011", 
						"00000001" when "00011100", 
						"00011111" when "00011101", 
						"00111101" when "00011110", 
						"00100011" when "00011111", 
						"01111011" when "00100000", 
						"01100101" when "00100001", 
						"01000111" when "00100010", 
						"01011001" when "00100011", 
						"00000011" when "00100100", 
						"00011101" when "00100101", 
						"00111111" when "00100110", 
						"00100001" when "00100111", 
						"10001011" when "00101000", 
						"10010101" when "00101001", 
						"10110111" when "00101010", 
						"10101001" when "00101011", 
						"11110011" when "00101100", 
						"11101101" when "00101101", 
						"11001111" when "00101110", 
						"11010001" when "00101111", 
						"11110010" when "00110000", 
						"11101100" when "00110001", 
						"11001110" when "00110010", 
						"11010000" when "00110011", 
						"10001010" when "00110100", 
						"10010100" when "00110101", 
						"10110110" when "00110110", 
						"10101000" when "00110111", 
						"00000010" when "00111000", 
						"00011100" when "00111001", 
						"00111110" when "00111010", 
						"00100000" when "00111011", 
						"01111010" when "00111100", 
						"01100100" when "00111101", 
						"01000110" when "00111110", 
						"01011000" when "00111111", 
						"11110110" when "01000000", 
						"11101000" when "01000001", 
						"11001010" when "01000010", 
						"11010100" when "01000011", 
						"10001110" when "01000100", 
						"10010000" when "01000101", 
						"10110010" when "01000110", 
						"10101100" when "01000111", 
						"00000110" when "01001000", 
						"00011000" when "01001001", 
						"00111010" when "01001010", 
						"00100100" when "01001011", 
						"01111110" when "01001100", 
						"01100000" when "01001101", 
						"01000010" when "01001110", 
						"01011100" when "01001111", 
						"01111111" when "01010000", 
						"01100001" when "01010001", 
						"01000011" when "01010010", 
						"01011101" when "01010011", 
						"00000111" when "01010100", 
						"00011001" when "01010101", 
						"00111011" when "01010110", 
						"00100101" when "01010111", 
						"10001111" when "01011000", 
						"10010001" when "01011001", 
						"10110011" when "01011010", 
						"10101101" when "01011011", 
						"11110111" when "01011100", 
						"11101001" when "01011101", 
						"11001011" when "01011110", 
						"11010101" when "01011111", 
						"10001101" when "01100000", 
						"10010011" when "01100001", 
						"10110001" when "01100010", 
						"10101111" when "01100011", 
						"11110101" when "01100100", 
						"11101011" when "01100101", 
						"11001001" when "01100110", 
						"11010111" when "01100111", 
						"01111101" when "01101000", 
						"01100011" when "01101001", 
						"01000001" when "01101010", 
						"01011111" when "01101011", 
						"00000101" when "01101100", 
						"00011011" when "01101101", 
						"00111001" when "01101110", 
						"00100111" when "01101111", 
						"00000100" when "01110000", 
						"00011010" when "01110001", 
						"00111000" when "01110010", 
						"00100110" when "01110011", 
						"01111100" when "01110100", 
						"01100010" when "01110101", 
						"01000000" when "01110110", 
						"01011110" when "01110111", 
						"11110100" when "01111000", 
						"11101010" when "01111001", 
						"11001000" when "01111010", 
						"11010110" when "01111011", 
						"10001100" when "01111100", 
						"10010010" when "01111101", 
						"10110000" when "01111110", 
						"10101110" when "01111111", 
						"10000101" when "10000000", 
						"10011011" when "10000001", 
						"10111001" when "10000010", 
						"10100111" when "10000011", 
						"11111101" when "10000100", 
						"11100011" when "10000101", 
						"11000001" when "10000110", 
						"11011111" when "10000111", 
						"01110101" when "10001000", 
						"01101011" when "10001001", 
						"01001001" when "10001010", 
						"01010111" when "10001011", 
						"00001101" when "10001100", 
						"00010011" when "10001101", 
						"00110001" when "10001110", 
						"00101111" when "10001111", 
						"00001100" when "10010000", 
						"00010010" when "10010001", 
						"00110000" when "10010010", 
						"00101110" when "10010011", 
						"01110100" when "10010100", 
						"01101010" when "10010101", 
						"01001000" when "10010110", 
						"01010110" when "10010111", 
						"11111100" when "10011000", 
						"11100010" when "10011001", 
						"11000000" when "10011010", 
						"11011110" when "10011011", 
						"10000100" when "10011100", 
						"10011010" when "10011101", 
						"10111000" when "10011110", 
						"10100110" when "10011111", 
						"11111110" when "10100000", 
						"11100000" when "10100001", 
						"11000010" when "10100010", 
						"11011100" when "10100011", 
						"10000110" when "10100100", 
						"10011000" when "10100101", 
						"10111010" when "10100110", 
						"10100100" when "10100111", 
						"00001110" when "10101000", 
						"00010000" when "10101001", 
						"00110010" when "10101010", 
						"00101100" when "10101011", 
						"01110110" when "10101100", 
						"01101000" when "10101101", 
						"01001010" when "10101110", 
						"01010100" when "10101111", 
						"01110111" when "10110000", 
						"01101001" when "10110001", 
						"01001011" when "10110010", 
						"01010101" when "10110011", 
						"00001111" when "10110100", 
						"00010001" when "10110101", 
						"00110011" when "10110110", 
						"00101101" when "10110111", 
						"10000111" when "10111000", 
						"10011001" when "10111001", 
						"10111011" when "10111010", 
						"10100101" when "10111011", 
						"11111111" when "10111100", 
						"11100001" when "10111101", 
						"11000011" when "10111110", 
						"11011101" when "10111111", 
						"01110011" when "11000000", 
						"01101101" when "11000001", 
						"01001111" when "11000010", 
						"01010001" when "11000011", 
						"00001011" when "11000100", 
						"00010101" when "11000101", 
						"00110111" when "11000110", 
						"00101001" when "11000111", 
						"10000011" when "11001000", 
						"10011101" when "11001001", 
						"10111111" when "11001010", 
						"10100001" when "11001011", 
						"11111011" when "11001100", 
						"11100101" when "11001101", 
						"11000111" when "11001110", 
						"11011001" when "11001111", 
						"11111010" when "11010000", 
						"11100100" when "11010001", 
						"11000110" when "11010010", 
						"11011000" when "11010011", 
						"10000010" when "11010100", 
						"10011100" when "11010101", 
						"10111110" when "11010110", 
						"10100000" when "11010111", 
						"00001010" when "11011000", 
						"00010100" when "11011001", 
						"00110110" when "11011010", 
						"00101000" when "11011011", 
						"01110010" when "11011100", 
						"01101100" when "11011101", 
						"01001110" when "11011110", 
						"01010000" when "11011111", 
						"00001000" when "11100000", 
						"00010110" when "11100001", 
						"00110100" when "11100010", 
						"00101010" when "11100011", 
						"01110000" when "11100100", 
						"01101110" when "11100101", 
						"01001100" when "11100110", 
						"01010010" when "11100111", 
						"11111000" when "11101000", 
						"11100110" when "11101001", 
						"11000100" when "11101010", 
						"11011010" when "11101011", 
						"10000000" when "11101100", 
						"10011110" when "11101101", 
						"10111100" when "11101110", 
						"10100010" when "11101111", 
						"10000001" when "11110000", 
						"10011111" when "11110001", 
						"10111101" when "11110010", 
						"10100011" when "11110011", 
						"11111001" when "11110100", 
						"11100111" when "11110101", 
						"11000101" when "11110110", 
						"11011011" when "11110111", 
						"01110001" when "11111000", 
						"01101111" when "11111001", 
						"01001101" when "11111010", 
						"01010011" when "11111011", 
						"00001001" when "11111100", 
						"00010111" when "11111101", 
						"00110101" when "11111110", 
						"00101011" when "11111111";

end mul_1E_mem;

