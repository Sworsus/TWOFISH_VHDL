----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:48:29 04/24/2021 
-- Design Name: 
-- Module Name:    mul_C6_mem - mul_C6_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_C6_mem is
	port (
			in_C6 : in STD_LOGIC_VECTOR (7 downto 0);
			out_C6 : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_C6_mem;

architecture mul_C6_mem of mul_C6_mem is

begin

	with in_C6 select
	out_C6 <= "00000000" when "00000000", 
				"11000110" when "00000001", 
				"11100101" when "00000010", 
				"00100011" when "00000011", 
				"10100011" when "00000100", 
				"01100101" when "00000101", 
				"01000110" when "00000110", 
				"10000000" when "00000111", 
				"00101111" when "00001000", 
				"11101001" when "00001001", 
				"11001010" when "00001010", 
				"00001100" when "00001011", 
				"10001100" when "00001100", 
				"01001010" when "00001101", 
				"01101001" when "00001110", 
				"10101111" when "00001111", 
				"01011110" when "00010000", 
				"10011000" when "00010001", 
				"10111011" when "00010010", 
				"01111101" when "00010011", 
				"11111101" when "00010100", 
				"00111011" when "00010101", 
				"00011000" when "00010110", 
				"11011110" when "00010111", 
				"01110001" when "00011000", 
				"10110111" when "00011001", 
				"10010100" when "00011010", 
				"01010010" when "00011011", 
				"11010010" when "00011100", 
				"00010100" when "00011101", 
				"00110111" when "00011110", 
				"11110001" when "00011111", 
				"10111100" when "00100000", 
				"01111010" when "00100001", 
				"01011001" when "00100010", 
				"10011111" when "00100011", 
				"00011111" when "00100100", 
				"11011001" when "00100101", 
				"11111010" when "00100110", 
				"00111100" when "00100111", 
				"10010011" when "00101000", 
				"01010101" when "00101001", 
				"01110110" when "00101010", 
				"10110000" when "00101011", 
				"00110000" when "00101100", 
				"11110110" when "00101101", 
				"11010101" when "00101110", 
				"00010011" when "00101111", 
				"11100010" when "00110000", 
				"00100100" when "00110001", 
				"00000111" when "00110010", 
				"11000001" when "00110011", 
				"01000001" when "00110100", 
				"10000111" when "00110101", 
				"10100100" when "00110110", 
				"01100010" when "00110111", 
				"11001101" when "00111000", 
				"00001011" when "00111001", 
				"00101000" when "00111010", 
				"11101110" when "00111011", 
				"01101110" when "00111100", 
				"10101000" when "00111101", 
				"10001011" when "00111110", 
				"01001101" when "00111111", 
				"00010001" when "01000000", 
				"11010111" when "01000001", 
				"11110100" when "01000010", 
				"00110010" when "01000011", 
				"10110010" when "01000100", 
				"01110100" when "01000101", 
				"01010111" when "01000110", 
				"10010001" when "01000111", 
				"00111110" when "01001000", 
				"11111000" when "01001001", 
				"11011011" when "01001010", 
				"00011101" when "01001011", 
				"10011101" when "01001100", 
				"01011011" when "01001101", 
				"01111000" when "01001110", 
				"10111110" when "01001111", 
				"01001111" when "01010000", 
				"10001001" when "01010001", 
				"10101010" when "01010010", 
				"01101100" when "01010011", 
				"11101100" when "01010100", 
				"00101010" when "01010101", 
				"00001001" when "01010110", 
				"11001111" when "01010111", 
				"01100000" when "01011000", 
				"10100110" when "01011001", 
				"10000101" when "01011010", 
				"01000011" when "01011011", 
				"11000011" when "01011100", 
				"00000101" when "01011101", 
				"00100110" when "01011110", 
				"11100000" when "01011111", 
				"10101101" when "01100000", 
				"01101011" when "01100001", 
				"01001000" when "01100010", 
				"10001110" when "01100011", 
				"00001110" when "01100100", 
				"11001000" when "01100101", 
				"11101011" when "01100110", 
				"00101101" when "01100111", 
				"10000010" when "01101000", 
				"01000100" when "01101001", 
				"01100111" when "01101010", 
				"10100001" when "01101011", 
				"00100001" when "01101100", 
				"11100111" when "01101101", 
				"11000100" when "01101110", 
				"00000010" when "01101111", 
				"11110011" when "01110000", 
				"00110101" when "01110001", 
				"00010110" when "01110010", 
				"11010000" when "01110011", 
				"01010000" when "01110100", 
				"10010110" when "01110101", 
				"10110101" when "01110110", 
				"01110011" when "01110111", 
				"11011100" when "01111000", 
				"00011010" when "01111001", 
				"00111001" when "01111010", 
				"11111111" when "01111011", 
				"01111111" when "01111100", 
				"10111001" when "01111101", 
				"10011010" when "01111110", 
				"01011100" when "01111111", 
				"00100010" when "10000000", 
				"11100100" when "10000001", 
				"11000111" when "10000010", 
				"00000001" when "10000011", 
				"10000001" when "10000100", 
				"01000111" when "10000101", 
				"01100100" when "10000110", 
				"10100010" when "10000111", 
				"00001101" when "10001000", 
				"11001011" when "10001001", 
				"11101000" when "10001010", 
				"00101110" when "10001011", 
				"10101110" when "10001100", 
				"01101000" when "10001101", 
				"01001011" when "10001110", 
				"10001101" when "10001111", 
				"01111100" when "10010000", 
				"10111010" when "10010001", 
				"10011001" when "10010010", 
				"01011111" when "10010011", 
				"11011111" when "10010100", 
				"00011001" when "10010101", 
				"00111010" when "10010110", 
				"11111100" when "10010111", 
				"01010011" when "10011000", 
				"10010101" when "10011001", 
				"10110110" when "10011010", 
				"01110000" when "10011011", 
				"11110000" when "10011100", 
				"00110110" when "10011101", 
				"00010101" when "10011110", 
				"11010011" when "10011111", 
				"10011110" when "10100000", 
				"01011000" when "10100001", 
				"01111011" when "10100010", 
				"10111101" when "10100011", 
				"00111101" when "10100100", 
				"11111011" when "10100101", 
				"11011000" when "10100110", 
				"00011110" when "10100111", 
				"10110001" when "10101000", 
				"01110111" when "10101001", 
				"01010100" when "10101010", 
				"10010010" when "10101011", 
				"00010010" when "10101100", 
				"11010100" when "10101101", 
				"11110111" when "10101110", 
				"00110001" when "10101111", 
				"11000000" when "10110000", 
				"00000110" when "10110001", 
				"00100101" when "10110010", 
				"11100011" when "10110011", 
				"01100011" when "10110100", 
				"10100101" when "10110101", 
				"10000110" when "10110110", 
				"01000000" when "10110111", 
				"11101111" when "10111000", 
				"00101001" when "10111001", 
				"00001010" when "10111010", 
				"11001100" when "10111011", 
				"01001100" when "10111100", 
				"10001010" when "10111101", 
				"10101001" when "10111110", 
				"01101111" when "10111111", 
				"00110011" when "11000000", 
				"11110101" when "11000001", 
				"11010110" when "11000010", 
				"00010000" when "11000011", 
				"10010000" when "11000100", 
				"01010110" when "11000101", 
				"01110101" when "11000110", 
				"10110011" when "11000111", 
				"00011100" when "11001000", 
				"11011010" when "11001001", 
				"11111001" when "11001010", 
				"00111111" when "11001011", 
				"10111111" when "11001100", 
				"01111001" when "11001101", 
				"01011010" when "11001110", 
				"10011100" when "11001111", 
				"01101101" when "11010000", 
				"10101011" when "11010001", 
				"10001000" when "11010010", 
				"01001110" when "11010011", 
				"11001110" when "11010100", 
				"00001000" when "11010101", 
				"00101011" when "11010110", 
				"11101101" when "11010111", 
				"01000010" when "11011000", 
				"10000100" when "11011001", 
				"10100111" when "11011010", 
				"01100001" when "11011011", 
				"11100001" when "11011100", 
				"00100111" when "11011101", 
				"00000100" when "11011110", 
				"11000010" when "11011111", 
				"10001111" when "11100000", 
				"01001001" when "11100001", 
				"01101010" when "11100010", 
				"10101100" when "11100011", 
				"00101100" when "11100100", 
				"11101010" when "11100101", 
				"11001001" when "11100110", 
				"00001111" when "11100111", 
				"10100000" when "11101000", 
				"01100110" when "11101001", 
				"01000101" when "11101010", 
				"10000011" when "11101011", 
				"00000011" when "11101100", 
				"11000101" when "11101101", 
				"11100110" when "11101110", 
				"00100000" when "11101111", 
				"11010001" when "11110000", 
				"00010111" when "11110001", 
				"00110100" when "11110010", 
				"11110010" when "11110011", 
				"01110010" when "11110100", 
				"10110100" when "11110101", 
				"10010111" when "11110110", 
				"01010001" when "11110111", 
				"11111110" when "11111000", 
				"00111000" when "11111001", 
				"00011011" when "11111010", 
				"11011101" when "11111011", 
				"01011101" when "11111100", 
				"10011011" when "11111101", 
				"10111000" when "11111110", 
				"01111110" when "11111111";

end mul_C6_mem;

