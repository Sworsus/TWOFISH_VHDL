----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:02:57 04/23/2021 
-- Design Name: 
-- Module Name:    mul_19_mem - mul_19_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_19_mem is
	port (
			in_19 : in STD_LOGIC_VECTOR (7 downto 0);
			out_19 : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_19_mem;

architecture mul_19_mem of mul_19_mem is

begin

	with in_19 select
		out_19 <= "00000000" when "00000000", "00011001" when "00000001", "00110010" when "00000010", "00101011" when "00000011",
					"01100100" when "00000100", "01111101" when "00000101", "01010110" when "00000110", "01001111" when "00000111",
					"11001000" when "00001000", "11010001" when "00001001", "11111010" when "00001010", "11100011" when "00001011",
					"10101100" when "00001100", "10110101" when "00001101", "10011110" when "00001110", "10000111" when "00001111",
					"11111001" when "00010000", "11100000" when "00010001", "11001011" when "00010010", "11010010" when "00010011",
					"10011101" when "00010100", "10000100" when "00010101", "10101111" when "00010110", "10110110" when "00010111",
					"00110001" when "00011000", "00101000" when "00011001", "00000011" when "00011010", "00011010" when "00011011",
					"01010101" when "00011100", "01001100" when "00011101", "01100111" when "00011110", "01111110" when "00011111",
					"10011011" when "00100000", "10000010" when "00100001", "10101001" when "00100010", "10110000" when "00100011",
					"11111111" when "00100100", "11100110" when "00100101", "11001101" when "00100110", "11010100" when "00100111",
					"01010011" when "00101000", "01001010" when "00101001", "01100001" when "00101010", "01111000" when "00101011",
					"00110111" when "00101100", "00101110" when "00101101", "00000101" when "00101110", "00011100" when "00101111",
					"01100010" when "00110000", "01111011" when "00110001", "01010000" when "00110010", "01001001" when "00110011",
					"00000110" when "00110100", "00011111" when "00110101", "00110100" when "00110110", "00101101" when "00110111",
					"10101010" when "00111000", "10110011" when "00111001", "10011000" when "00111010", "10000001" when "00111011",
					"11001110" when "00111100", "11010111" when "00111101", "11111100" when "00111110", "11100101" when "00111111",
					"01011111" when "01000000", "01000110" when "01000001", "01101101" when "01000010", "01110100" when "01000011",
					"00111011" when "01000100", "00100010" when "01000101", "00001001" when "01000110", "00010000" when "01000111",
					"10010111" when "01001000", "10001110" when "01001001", "10100101" when "01001010", "10111100" when "01001011",
					"11110011" when "01001100", "11101010" when "01001101", "11000001" when "01001110", "11011000" when "01001111",
					"10100110" when "01010000", "10111111" when "01010001", "10010100" when "01010010", "10001101" when "01010011",
					"11000010" when "01010100", "11011011" when "01010101", "11110000" when "01010110", "11101001" when "01010111",
					"01101110" when "01011000", "01110111" when "01011001", "01011100" when "01011010", "01000101" when "01011011",
					"00001010" when "01011100", "00010011" when "01011101", "00111000" when "01011110", "00100001" when "01011111",
					"11000100" when "01100000", "11011101" when "01100001", "11110110" when "01100010", "11101111" when "01100011",
					"10100000" when "01100100", "10111001" when "01100101", "10010010" when "01100110", "10001011" when "01100111",
					"00001100" when "01101000", "00010101" when "01101001", "00111110" when "01101010", "00100111" when "01101011",
					"01101000" when "01101100", "01110001" when "01101101", "01011010" when "01101110", "01000011" when "01101111",
					"00111101" when "01110000", "00100100" when "01110001", "00001111" when "01110010", "00010110" when "01110011",
					"01011001" when "01110100", "01000000" when "01110101", "01101011" when "01110110", "01110010" when "01110111",
					"11110101" when "01111000", "11101100" when "01111001", "11000111" when "01111010", "11011110" when "01111011",
					"10010001" when "01111100", "10001000" when "01111101", "10100011" when "01111110", "10111010" when "01111111",
					"10111110" when "10000000", "10100111" when "10000001", "10001100" when "10000010", "10010101" when "10000011",
					"11011010" when "10000100", "11000011" when "10000101", "11101000" when "10000110", "11110001" when "10000111",
					"01110110" when "10001000", "01101111" when "10001001", "01000100" when "10001010", "01011101" when "10001011",
					"00010010" when "10001100", "00001011" when "10001101", "00100000" when "10001110", "00111001" when "10001111",
					"01000111" when "10010000", "01011110" when "10010001", "01110101" when "10010010", "01101100" when "10010011",
					"00100011" when "10010100", "00111010" when "10010101", "00010001" when "10010110", "00001000" when "10010111",
					"10001111" when "10011000", "10010110" when "10011001", "10111101" when "10011010", "10100100" when "10011011",
					"11101011" when "10011100", "11110010" when "10011101", "11011001" when "10011110", "11000000" when "10011111",
					"00100101" when "10100000", "00111100" when "10100001", "00010111" when "10100010", "00001110" when "10100011",
					"01000001" when "10100100", "01011000" when "10100101", "01110011" when "10100110", "01101010" when "10100111",
					"11101101" when "10101000", "11110100" when "10101001", "11011111" when "10101010", "11000110" when "10101011",
					"10001001" when "10101100", "10010000" when "10101101", "10111011" when "10101110", "10100010" when "10101111",
					"11011100" when "10110000", "11000101" when "10110001", "11101110" when "10110010", "11110111" when "10110011",
					"10111000" when "10110100", "10100001" when "10110101", "10001010" when "10110110", "10010011" when "10110111",
					"00010100" when "10111000", "00001101" when "10111001", "00100110" when "10111010", "00111111" when "10111011",
					"01110000" when "10111100", "01101001" when "10111101", "01000010" when "10111110", "01011011" when "10111111",
					"11100001" when "11000000", "11111000" when "11000001", "11010011" when "11000010", "11001010" when "11000011",
					"10000101" when "11000100", "10011100" when "11000101", "10110111" when "11000110", "10101110" when "11000111",
					"00101001" when "11001000", "00110000" when "11001001", "00011011" when "11001010", "00000010" when "11001011",
					"01001101" when "11001100", "01010100" when "11001101", "01111111" when "11001110", "01100110" when "11001111",
					"00011000" when "11010000", "00000001" when "11010001", "00101010" when "11010010", "00110011" when "11010011",
					"01111100" when "11010100", "01100101" when "11010101", "01001110" when "11010110", "01010111" when "11010111",
					"11010000" when "11011000", "11001001" when "11011001", "11100010" when "11011010", "11111011" when "11011011",
					"10110100" when "11011100", "10101101" when "11011101", "10000110" when "11011110", "10011111" when "11011111",
					"01111010" when "11100000", "01100011" when "11100001", "01001000" when "11100010", "01010001" when "11100011",
					"00011110" when "11100100", "00000111" when "11100101", "00101100" when "11100110", "00110101" when "11100111",
					"10110010" when "11101000", "10101011" when "11101001", "10000000" when "11101010", "10011001" when "11101011",
					"11010110" when "11101100", "11001111" when "11101101", "11100100" when "11101110", "11111101" when "11101111",
					"10000011" when "11110000", "10011010" when "11110001", "10110001" when "11110010", "10101000" when "11110011",
					"11100111" when "11110100", "11111110" when "11110101", "11010101" when "11110110", "11001100" when "11110111",
					"01001011" when "11111000", "01010010" when "11111001", "01111001" when "11111010", "01100000" when "11111011",
					"00101111" when "11111100", "00110110" when "11111101", "00011101" when "11111110", "00000100" when "11111111";

end mul_19_mem;

