----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    01:00:50 04/24/2021 
-- Design Name: 
-- Module Name:    mul_55_mem - mul_55_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity mul_55_mem is
	port (
			in_55 : in STD_LOGIC_VECTOR (7 downto 0);
			out_55 : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_55_mem;

architecture mul_55_mem of mul_55_mem is
begin

	with in_55 select
	out_55 <= "00000000" when "00000000", 
				"01010101" when "00000001", 
				"10101010" when "00000010", 
				"11111111" when "00000011", 
				"00111101" when "00000100", 
				"01101000" when "00000101", 
				"10010111" when "00000110", 
				"11000010" when "00000111", 
				"01111010" when "00001000", 
				"00101111" when "00001001", 
				"11010000" when "00001010", 
				"10000101" when "00001011", 
				"01000111" when "00001100", 
				"00010010" when "00001101", 
				"11101101" when "00001110", 
				"10111000" when "00001111", 
				"11110100" when "00010000", 
				"10100001" when "00010001", 
				"01011110" when "00010010", 
				"00001011" when "00010011", 
				"11001001" when "00010100", 
				"10011100" when "00010101", 
				"01100011" when "00010110", 
				"00110110" when "00010111", 
				"10001110" when "00011000", 
				"11011011" when "00011001", 
				"00100100" when "00011010", 
				"01110001" when "00011011", 
				"10110011" when "00011100", 
				"11100110" when "00011101", 
				"00011001" when "00011110", 
				"01001100" when "00011111", 
				"10000001" when "00100000", 
				"11010100" when "00100001", 
				"00101011" when "00100010", 
				"01111110" when "00100011", 
				"10111100" when "00100100", 
				"11101001" when "00100101", 
				"00010110" when "00100110", 
				"01000011" when "00100111", 
				"11111011" when "00101000", 
				"10101110" when "00101001", 
				"01010001" when "00101010", 
				"00000100" when "00101011", 
				"11000110" when "00101100", 
				"10010011" when "00101101", 
				"01101100" when "00101110", 
				"00111001" when "00101111", 
				"01110101" when "00110000", 
				"00100000" when "00110001", 
				"11011111" when "00110010", 
				"10001010" when "00110011", 
				"01001000" when "00110100", 
				"00011101" when "00110101", 
				"11100010" when "00110110", 
				"10110111" when "00110111", 
				"00001111" when "00111000", 
				"01011010" when "00111001", 
				"10100101" when "00111010", 
				"11110000" when "00111011", 
				"00110010" when "00111100", 
				"01100111" when "00111101", 
				"10011000" when "00111110", 
				"11001101" when "00111111", 
				"01101011" when "01000000", 
				"00111110" when "01000001", 
				"11000001" when "01000010", 
				"10010100" when "01000011", 
				"01010110" when "01000100", 
				"00000011" when "01000101", 
				"11111100" when "01000110", 
				"10101001" when "01000111", 
				"00010001" when "01001000", 
				"01000100" when "01001001", 
				"10111011" when "01001010", 
				"11101110" when "01001011", 
				"00101100" when "01001100", 
				"01111001" when "01001101", 
				"10000110" when "01001110", 
				"11010011" when "01001111", 
				"10011111" when "01010000", 
				"11001010" when "01010001", 
				"00110101" when "01010010", 
				"01100000" when "01010011", 
				"10100010" when "01010100", 
				"11110111" when "01010101", 
				"00001000" when "01010110", 
				"01011101" when "01010111", 
				"11100101" when "01011000", 
				"10110000" when "01011001", 
				"01001111" when "01011010", 
				"00011010" when "01011011", 
				"11011000" when "01011100", 
				"10001101" when "01011101", 
				"01110010" when "01011110", 
				"00100111" when "01011111", 
				"11101010" when "01100000", 
				"10111111" when "01100001", 
				"01000000" when "01100010", 
				"00010101" when "01100011", 
				"11010111" when "01100100", 
				"10000010" when "01100101", 
				"01111101" when "01100110", 
				"00101000" when "01100111", 
				"10010000" when "01101000", 
				"11000101" when "01101001", 
				"00111010" when "01101010", 
				"01101111" when "01101011", 
				"10101101" when "01101100", 
				"11111000" when "01101101", 
				"00000111" when "01101110", 
				"01010010" when "01101111", 
				"00011110" when "01110000", 
				"01001011" when "01110001", 
				"10110100" when "01110010", 
				"11100001" when "01110011", 
				"00100011" when "01110100", 
				"01110110" when "01110101", 
				"10001001" when "01110110", 
				"11011100" when "01110111", 
				"01100100" when "01111000", 
				"00110001" when "01111001", 
				"11001110" when "01111010", 
				"10011011" when "01111011", 
				"01011001" when "01111100", 
				"00001100" when "01111101", 
				"11110011" when "01111110", 
				"10100110" when "01111111", 
				"11010110" when "10000000", 
				"10000011" when "10000001", 
				"01111100" when "10000010", 
				"00101001" when "10000011", 
				"11101011" when "10000100", 
				"10111110" when "10000101", 
				"01000001" when "10000110", 
				"00010100" when "10000111", 
				"10101100" when "10001000", 
				"11111001" when "10001001", 
				"00000110" when "10001010", 
				"01010011" when "10001011", 
				"10010001" when "10001100", 
				"11000100" when "10001101", 
				"00111011" when "10001110", 
				"01101110" when "10001111", 
				"00100010" when "10010000", 
				"01110111" when "10010001", 
				"10001000" when "10010010", 
				"11011101" when "10010011", 
				"00011111" when "10010100", 
				"01001010" when "10010101", 
				"10110101" when "10010110", 
				"11100000" when "10010111", 
				"01011000" when "10011000", 
				"00001101" when "10011001", 
				"11110010" when "10011010", 
				"10100111" when "10011011", 
				"01100101" when "10011100", 
				"00110000" when "10011101", 
				"11001111" when "10011110", 
				"10011010" when "10011111", 
				"01010111" when "10100000", 
				"00000010" when "10100001", 
				"11111101" when "10100010", 
				"10101000" when "10100011", 
				"01101010" when "10100100", 
				"00111111" when "10100101", 
				"11000000" when "10100110", 
				"10010101" when "10100111", 
				"00101101" when "10101000", 
				"01111000" when "10101001", 
				"10000111" when "10101010", 
				"11010010" when "10101011", 
				"00010000" when "10101100", 
				"01000101" when "10101101", 
				"10111010" when "10101110", 
				"11101111" when "10101111", 
				"10100011" when "10110000", 
				"11110110" when "10110001", 
				"00001001" when "10110010", 
				"01011100" when "10110011", 
				"10011110" when "10110100", 
				"11001011" when "10110101", 
				"00110100" when "10110110", 
				"01100001" when "10110111", 
				"11011001" when "10111000", 
				"10001100" when "10111001", 
				"01110011" when "10111010", 
				"00100110" when "10111011", 
				"11100100" when "10111100", 
				"10110001" when "10111101", 
				"01001110" when "10111110", 
				"00011011" when "10111111", 
				"10111101" when "11000000", 
				"11101000" when "11000001", 
				"00010111" when "11000010", 
				"01000010" when "11000011", 
				"10000000" when "11000100", 
				"11010101" when "11000101", 
				"00101010" when "11000110", 
				"01111111" when "11000111", 
				"11000111" when "11001000", 
				"10010010" when "11001001", 
				"01101101" when "11001010", 
				"00111000" when "11001011", 
				"11111010" when "11001100", 
				"10101111" when "11001101", 
				"01010000" when "11001110", 
				"00000101" when "11001111", 
				"01001001" when "11010000", 
				"00011100" when "11010001", 
				"11100011" when "11010010", 
				"10110110" when "11010011", 
				"01110100" when "11010100", 
				"00100001" when "11010101", 
				"11011110" when "11010110", 
				"10001011" when "11010111", 
				"00110011" when "11011000", 
				"01100110" when "11011001", 
				"10011001" when "11011010", 
				"11001100" when "11011011", 
				"00001110" when "11011100", 
				"01011011" when "11011101", 
				"10100100" when "11011110", 
				"11110001" when "11011111", 
				"00111100" when "11100000", 
				"01101001" when "11100001", 
				"10010110" when "11100010", 
				"11000011" when "11100011", 
				"00000001" when "11100100", 
				"01010100" when "11100101", 
				"10101011" when "11100110", 
				"11111110" when "11100111", 
				"01000110" when "11101000", 
				"00010011" when "11101001", 
				"11101100" when "11101010", 
				"10111001" when "11101011", 
				"01111011" when "11101100", 
				"00101110" when "11101101", 
				"11010001" when "11101110", 
				"10000100" when "11101111", 
				"11001000" when "11110000", 
				"10011101" when "11110001", 
				"01100010" when "11110010", 
				"00110111" when "11110011", 
				"11110101" when "11110100", 
				"10100000" when "11110101", 
				"01011111" when "11110110", 
				"00001010" when "11110111", 
				"10110010" when "11111000", 
				"11100111" when "11111001", 
				"00011000" when "11111010", 
				"01001101" when "11111011", 
				"10001111" when "11111100", 
				"11011010" when "11111101", 
				"00100101" when "11111110", 
				"01110000" when "11111111";

end mul_55_mem;

