----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    01:32:05 04/24/2021 
-- Design Name: 
-- Module Name:    mul_58_mem - mul_58_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_58_mem is
	port (
			in_58 : in STD_LOGIC_VECTOR (7 downto 0);
			out_58 : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_58_mem;

architecture mul_58_mem of mul_58_mem is

begin

	with in_58 select
	out_58 <= "00000000" when "00000000", 
				"01011000" when "00000001", 
				"10110000" when "00000010", 
				"11101000" when "00000011", 
				"00001001" when "00000100", 
				"01010001" when "00000101", 
				"10111001" when "00000110", 
				"11100001" when "00000111", 
				"00010010" when "00001000", 
				"01001010" when "00001001", 
				"10100010" when "00001010", 
				"11111010" when "00001011", 
				"00011011" when "00001100", 
				"01000011" when "00001101", 
				"10101011" when "00001110", 
				"11110011" when "00001111", 
				"00100100" when "00010000", 
				"01111100" when "00010001", 
				"10010100" when "00010010", 
				"11001100" when "00010011", 
				"00101101" when "00010100", 
				"01110101" when "00010101", 
				"10011101" when "00010110", 
				"11000101" when "00010111", 
				"00110110" when "00011000", 
				"01101110" when "00011001", 
				"10000110" when "00011010", 
				"11011110" when "00011011", 
				"00111111" when "00011100", 
				"01100111" when "00011101", 
				"10001111" when "00011110", 
				"11010111" when "00011111", 
				"01001000" when "00100000", 
				"00010000" when "00100001", 
				"11111000" when "00100010", 
				"10100000" when "00100011", 
				"01000001" when "00100100", 
				"00011001" when "00100101", 
				"11110001" when "00100110", 
				"10101001" when "00100111", 
				"01011010" when "00101000", 
				"00000010" when "00101001", 
				"11101010" when "00101010", 
				"10110010" when "00101011", 
				"01010011" when "00101100", 
				"00001011" when "00101101", 
				"11100011" when "00101110", 
				"10111011" when "00101111", 
				"01101100" when "00110000", 
				"00110100" when "00110001", 
				"11011100" when "00110010", 
				"10000100" when "00110011", 
				"01100101" when "00110100", 
				"00111101" when "00110101", 
				"11010101" when "00110110", 
				"10001101" when "00110111", 
				"01111110" when "00111000", 
				"00100110" when "00111001", 
				"11001110" when "00111010", 
				"10010110" when "00111011", 
				"01110111" when "00111100", 
				"00101111" when "00111101", 
				"11000111" when "00111110", 
				"10011111" when "00111111", 
				"10010000" when "01000000", 
				"11001000" when "01000001", 
				"00100000" when "01000010", 
				"01111000" when "01000011", 
				"10011001" when "01000100", 
				"11000001" when "01000101", 
				"00101001" when "01000110", 
				"01110001" when "01000111", 
				"10000010" when "01001000", 
				"11011010" when "01001001", 
				"00110010" when "01001010", 
				"01101010" when "01001011", 
				"10001011" when "01001100", 
				"11010011" when "01001101", 
				"00111011" when "01001110", 
				"01100011" when "01001111", 
				"10110100" when "01010000", 
				"11101100" when "01010001", 
				"00000100" when "01010010", 
				"01011100" when "01010011", 
				"10111101" when "01010100", 
				"11100101" when "01010101", 
				"00001101" when "01010110", 
				"01010101" when "01010111", 
				"10100110" when "01011000", 
				"11111110" when "01011001", 
				"00010110" when "01011010", 
				"01001110" when "01011011", 
				"10101111" when "01011100", 
				"11110111" when "01011101", 
				"00011111" when "01011110", 
				"01000111" when "01011111", 
				"11011000" when "01100000", 
				"10000000" when "01100001", 
				"01101000" when "01100010", 
				"00110000" when "01100011", 
				"11010001" when "01100100", 
				"10001001" when "01100101", 
				"01100001" when "01100110", 
				"00111001" when "01100111", 
				"11001010" when "01101000", 
				"10010010" when "01101001", 
				"01111010" when "01101010", 
				"00100010" when "01101011", 
				"11000011" when "01101100", 
				"10011011" when "01101101", 
				"01110011" when "01101110", 
				"00101011" when "01101111", 
				"11111100" when "01110000", 
				"10100100" when "01110001", 
				"01001100" when "01110010", 
				"00010100" when "01110011", 
				"11110101" when "01110100", 
				"10101101" when "01110101", 
				"01000101" when "01110110", 
				"00011101" when "01110111", 
				"11101110" when "01111000", 
				"10110110" when "01111001", 
				"01011110" when "01111010", 
				"00000110" when "01111011", 
				"11100111" when "01111100", 
				"10111111" when "01111101", 
				"01010111" when "01111110", 
				"00001111" when "01111111", 
				"01001001" when "10000000", 
				"00010001" when "10000001", 
				"11111001" when "10000010", 
				"10100001" when "10000011", 
				"01000000" when "10000100", 
				"00011000" when "10000101", 
				"11110000" when "10000110", 
				"10101000" when "10000111", 
				"01011011" when "10001000", 
				"00000011" when "10001001", 
				"11101011" when "10001010", 
				"10110011" when "10001011", 
				"01010010" when "10001100", 
				"00001010" when "10001101", 
				"11100010" when "10001110", 
				"10111010" when "10001111", 
				"01101101" when "10010000", 
				"00110101" when "10010001", 
				"11011101" when "10010010", 
				"10000101" when "10010011", 
				"01100100" when "10010100", 
				"00111100" when "10010101", 
				"11010100" when "10010110", 
				"10001100" when "10010111", 
				"01111111" when "10011000", 
				"00100111" when "10011001", 
				"11001111" when "10011010", 
				"10010111" when "10011011", 
				"01110110" when "10011100", 
				"00101110" when "10011101", 
				"11000110" when "10011110", 
				"10011110" when "10011111", 
				"00000001" when "10100000", 
				"01011001" when "10100001", 
				"10110001" when "10100010", 
				"11101001" when "10100011", 
				"00001000" when "10100100", 
				"01010000" when "10100101", 
				"10111000" when "10100110", 
				"11100000" when "10100111", 
				"00010011" when "10101000", 
				"01001011" when "10101001", 
				"10100011" when "10101010", 
				"11111011" when "10101011", 
				"00011010" when "10101100", 
				"01000010" when "10101101", 
				"10101010" when "10101110", 
				"11110010" when "10101111", 
				"00100101" when "10110000", 
				"01111101" when "10110001", 
				"10010101" when "10110010", 
				"11001101" when "10110011", 
				"00101100" when "10110100", 
				"01110100" when "10110101", 
				"10011100" when "10110110", 
				"11000100" when "10110111", 
				"00110111" when "10111000", 
				"01101111" when "10111001", 
				"10000111" when "10111010", 
				"11011111" when "10111011", 
				"00111110" when "10111100", 
				"01100110" when "10111101", 
				"10001110" when "10111110", 
				"11010110" when "10111111", 
				"11011001" when "11000000", 
				"10000001" when "11000001", 
				"01101001" when "11000010", 
				"00110001" when "11000011", 
				"11010000" when "11000100", 
				"10001000" when "11000101", 
				"01100000" when "11000110", 
				"00111000" when "11000111", 
				"11001011" when "11001000", 
				"10010011" when "11001001", 
				"01111011" when "11001010", 
				"00100011" when "11001011", 
				"11000010" when "11001100", 
				"10011010" when "11001101", 
				"01110010" when "11001110", 
				"00101010" when "11001111", 
				"11111101" when "11010000", 
				"10100101" when "11010001", 
				"01001101" when "11010010", 
				"00010101" when "11010011", 
				"11110100" when "11010100", 
				"10101100" when "11010101", 
				"01000100" when "11010110", 
				"00011100" when "11010111", 
				"11101111" when "11011000", 
				"10110111" when "11011001", 
				"01011111" when "11011010", 
				"00000111" when "11011011", 
				"11100110" when "11011100", 
				"10111110" when "11011101", 
				"01010110" when "11011110", 
				"00001110" when "11011111", 
				"10010001" when "11100000", 
				"11001001" when "11100001", 
				"00100001" when "11100010", 
				"01111001" when "11100011", 
				"10011000" when "11100100", 
				"11000000" when "11100101", 
				"00101000" when "11100110", 
				"01110000" when "11100111", 
				"10000011" when "11101000", 
				"11011011" when "11101001", 
				"00110011" when "11101010", 
				"01101011" when "11101011", 
				"10001010" when "11101100", 
				"11010010" when "11101101", 
				"00111010" when "11101110", 
				"01100010" when "11101111", 
				"10110101" when "11110000", 
				"11101101" when "11110001", 
				"00000101" when "11110010", 
				"01011101" when "11110011", 
				"10111100" when "11110100", 
				"11100100" when "11110101", 
				"00001100" when "11110110", 
				"01010100" when "11110111", 
				"10100111" when "11111000", 
				"11111111" when "11111001", 
				"00010111" when "11111010", 
				"01001111" when "11111011", 
				"10101110" when "11111100", 
				"11110110" when "11111101", 
				"00011110" when "11111110", 
				"01000110" when "11111111";

end mul_58_mem;

