----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:15:56 04/24/2021 
-- Design Name: 
-- Module Name:    mul_A4_mem - mul_A4_mem 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mul_A4_mem is
	port (
			in_A4 : in STD_LOGIC_VECTOR (7 downto 0);
			out_A4 : out STD_LOGIC_VECTOR (7 downto 0)
			);
end mul_A4_mem;

architecture mul_A4_mem of mul_A4_mem is

begin

	with in_A4 select
	out_A4 <= "00000000" when "00000000", 
				"10100100" when "00000001", 
				"00100001" when "00000010", 
				"10000101" when "00000011", 
				"01000010" when "00000100", 
				"11100110" when "00000101", 
				"01100011" when "00000110", 
				"11000111" when "00000111", 
				"10000100" when "00001000", 
				"00100000" when "00001001", 
				"10100101" when "00001010", 
				"00000001" when "00001011", 
				"11000110" when "00001100", 
				"01100010" when "00001101", 
				"11100111" when "00001110", 
				"01000011" when "00001111", 
				"01100001" when "00010000", 
				"11000101" when "00010001", 
				"01000000" when "00010010", 
				"11100100" when "00010011", 
				"00100011" when "00010100", 
				"10000111" when "00010101", 
				"00000010" when "00010110", 
				"10100110" when "00010111", 
				"11100101" when "00011000", 
				"01000001" when "00011001", 
				"11000100" when "00011010", 
				"01100000" when "00011011", 
				"10100111" when "00011100", 
				"00000011" when "00011101", 
				"10000110" when "00011110", 
				"00100010" when "00011111", 
				"11000010" when "00100000", 
				"01100110" when "00100001", 
				"11100011" when "00100010", 
				"01000111" when "00100011", 
				"10000000" when "00100100", 
				"00100100" when "00100101", 
				"10100001" when "00100110", 
				"00000101" when "00100111", 
				"01000110" when "00101000", 
				"11100010" when "00101001", 
				"01100111" when "00101010", 
				"11000011" when "00101011", 
				"00000100" when "00101100", 
				"10100000" when "00101101", 
				"00100101" when "00101110", 
				"10000001" when "00101111", 
				"10100011" when "00110000", 
				"00000111" when "00110001", 
				"10000010" when "00110010", 
				"00100110" when "00110011", 
				"11100001" when "00110100", 
				"01000101" when "00110101", 
				"11000000" when "00110110", 
				"01100100" when "00110111", 
				"00100111" when "00111000", 
				"10000011" when "00111001", 
				"00000110" when "00111010", 
				"10100010" when "00111011", 
				"01100101" when "00111100", 
				"11000001" when "00111101", 
				"01000100" when "00111110", 
				"11100000" when "00111111", 
				"11101101" when "01000000", 
				"01001001" when "01000001", 
				"11001100" when "01000010", 
				"01101000" when "01000011", 
				"10101111" when "01000100", 
				"00001011" when "01000101", 
				"10001110" when "01000110", 
				"00101010" when "01000111", 
				"01101001" when "01001000", 
				"11001101" when "01001001", 
				"01001000" when "01001010", 
				"11101100" when "01001011", 
				"00101011" when "01001100", 
				"10001111" when "01001101", 
				"00001010" when "01001110", 
				"10101110" when "01001111", 
				"10001100" when "01010000", 
				"00101000" when "01010001", 
				"10101101" when "01010010", 
				"00001001" when "01010011", 
				"11001110" when "01010100", 
				"01101010" when "01010101", 
				"11101111" when "01010110", 
				"01001011" when "01010111", 
				"00001000" when "01011000", 
				"10101100" when "01011001", 
				"00101001" when "01011010", 
				"10001101" when "01011011", 
				"01001010" when "01011100", 
				"11101110" when "01011101", 
				"01101011" when "01011110", 
				"11001111" when "01011111", 
				"00101111" when "01100000", 
				"10001011" when "01100001", 
				"00001110" when "01100010", 
				"10101010" when "01100011", 
				"01101101" when "01100100", 
				"11001001" when "01100101", 
				"01001100" when "01100110", 
				"11101000" when "01100111", 
				"10101011" when "01101000", 
				"00001111" when "01101001", 
				"10001010" when "01101010", 
				"00101110" when "01101011", 
				"11101001" when "01101100", 
				"01001101" when "01101101", 
				"11001000" when "01101110", 
				"01101100" when "01101111", 
				"01001110" when "01110000", 
				"11101010" when "01110001", 
				"01101111" when "01110010", 
				"11001011" when "01110011", 
				"00001100" when "01110100", 
				"10101000" when "01110101", 
				"00101101" when "01110110", 
				"10001001" when "01110111", 
				"11001010" when "01111000", 
				"01101110" when "01111001", 
				"11101011" when "01111010", 
				"01001111" when "01111011", 
				"10001000" when "01111100", 
				"00101100" when "01111101", 
				"10101001" when "01111110", 
				"00001101" when "01111111", 
				"10110011" when "10000000", 
				"00010111" when "10000001", 
				"10010010" when "10000010", 
				"00110110" when "10000011", 
				"11110001" when "10000100", 
				"01010101" when "10000101", 
				"11010000" when "10000110", 
				"01110100" when "10000111", 
				"00110111" when "10001000", 
				"10010011" when "10001001", 
				"00010110" when "10001010", 
				"10110010" when "10001011", 
				"01110101" when "10001100", 
				"11010001" when "10001101", 
				"01010100" when "10001110", 
				"11110000" when "10001111", 
				"11010010" when "10010000", 
				"01110110" when "10010001", 
				"11110011" when "10010010", 
				"01010111" when "10010011", 
				"10010000" when "10010100", 
				"00110100" when "10010101", 
				"10110001" when "10010110", 
				"00010101" when "10010111", 
				"01010110" when "10011000", 
				"11110010" when "10011001", 
				"01110111" when "10011010", 
				"11010011" when "10011011", 
				"00010100" when "10011100", 
				"10110000" when "10011101", 
				"00110101" when "10011110", 
				"10010001" when "10011111", 
				"01110001" when "10100000", 
				"11010101" when "10100001", 
				"01010000" when "10100010", 
				"11110100" when "10100011", 
				"00110011" when "10100100", 
				"10010111" when "10100101", 
				"00010010" when "10100110", 
				"10110110" when "10100111", 
				"11110101" when "10101000", 
				"01010001" when "10101001", 
				"11010100" when "10101010", 
				"01110000" when "10101011", 
				"10110111" when "10101100", 
				"00010011" when "10101101", 
				"10010110" when "10101110", 
				"00110010" when "10101111", 
				"00010000" when "10110000", 
				"10110100" when "10110001", 
				"00110001" when "10110010", 
				"10010101" when "10110011", 
				"01010010" when "10110100", 
				"11110110" when "10110101", 
				"01110011" when "10110110", 
				"11010111" when "10110111", 
				"10010100" when "10111000", 
				"00110000" when "10111001", 
				"10110101" when "10111010", 
				"00010001" when "10111011", 
				"11010110" when "10111100", 
				"01110010" when "10111101", 
				"11110111" when "10111110", 
				"01010011" when "10111111", 
				"01011110" when "11000000", 
				"11111010" when "11000001", 
				"01111111" when "11000010", 
				"11011011" when "11000011", 
				"00011100" when "11000100", 
				"10111000" when "11000101", 
				"00111101" when "11000110", 
				"10011001" when "11000111", 
				"11011010" when "11001000", 
				"01111110" when "11001001", 
				"11111011" when "11001010", 
				"01011111" when "11001011", 
				"10011000" when "11001100", 
				"00111100" when "11001101", 
				"10111001" when "11001110", 
				"00011101" when "11001111", 
				"00111111" when "11010000", 
				"10011011" when "11010001", 
				"00011110" when "11010010", 
				"10111010" when "11010011", 
				"01111101" when "11010100", 
				"11011001" when "11010101", 
				"01011100" when "11010110", 
				"11111000" when "11010111", 
				"10111011" when "11011000", 
				"00011111" when "11011001", 
				"10011010" when "11011010", 
				"00111110" when "11011011", 
				"11111001" when "11011100", 
				"01011101" when "11011101", 
				"11011000" when "11011110", 
				"01111100" when "11011111", 
				"10011100" when "11100000", 
				"00111000" when "11100001", 
				"10111101" when "11100010", 
				"00011001" when "11100011", 
				"11011110" when "11100100", 
				"01111010" when "11100101", 
				"11111111" when "11100110", 
				"01011011" when "11100111", 
				"00011000" when "11101000", 
				"10111100" when "11101001", 
				"00111001" when "11101010", 
				"10011101" when "11101011", 
				"01011010" when "11101100", 
				"11111110" when "11101101", 
				"01111011" when "11101110", 
				"11011111" when "11101111", 
				"11111101" when "11110000", 
				"01011001" when "11110001", 
				"11011100" when "11110010", 
				"01111000" when "11110011", 
				"10111111" when "11110100", 
				"00011011" when "11110101", 
				"10011110" when "11110110", 
				"00111010" when "11110111", 
				"01111001" when "11111000", 
				"11011101" when "11111001", 
				"01011000" when "11111010", 
				"11111100" when "11111011", 
				"00111011" when "11111100", 
				"10011111" when "11111101", 
				"00011010" when "11111110", 
				"10111110" when "11111111";

end mul_A4_mem;

